module bit_stream (
    input clk,
    input EA,
    input [10:0] count_h,
    input [10:0] count_v,
    input [8:0] platform_const_h_0,
    input [8:0] platform_const_v_0,
    input [8:0] platform_const_h_1,
    input [8:0] platform_const_v_1,
    input [8:0] platform_const_h_2,
    input [8:0] platform_const_v_2,
    input [8:0] platform_const_h_3,
    input [8:0] platform_const_v_3,
    input [8:0] ground_h,
    input [8:0] ground_v,
    input [8:0] jump,
    input game_over,
    input [8:0] shift_h,
    input sprite_choice,
    output reg r, g, b
);

	// Registers to draw sprites
	reg doodle_sprite [0:1][0:80][0:80];
	reg platform_sprite [0:3][0:100][0:30];
	integer i = 0;
	reg [8:0] platform_v [0:3], platform_h[0:3];
	integer platform_const_v[0:3], platform_const_h[0:3];
	integer doodle_h, doodle_v;

	always @ (posedge clk)
	begin
			
			if (EA) begin
				if (!game_over) begin
					if (count_h >= 0) begin //background painting
						r = 1;
						g = 1;
						b = 1;
					end //---
						//setting doodle's coordinates:
					//horizontal: with constant shift & user's control shift
					//vertical: with jump & current platform vertical coordinates
					doodle_h = count_h - ground_h + shift_h - 600;
					doodle_v = count_v - ground_v - jump - 200;
					platform_const_v[0] = platform_const_v_0;
					platform_const_h[0] = platform_const_h_0;
							
					platform_const_v[1] = platform_const_v_1;
					platform_const_h[1] = platform_const_h_1;
							
					platform_const_v[2] = platform_const_v_2;
					platform_const_h[2] = platform_const_h_2;
							
					platform_const_v[3] = platform_const_v_3;
					platform_const_h[3] = platform_const_h_3;
					//setting platform coordinates with constant shifts
				for (i = 0; i < 4; i = i + 1) begin
					platform_h[i] = count_h - platform_const_h[i];
					platform_v[i] = count_v - platform_const_v[i];
					end	
					
					//assigning 1 to black pixels and 2 to green pixels inside of doodle
					doodle_sprite[0][4][16] = 2; doodle_sprite[0][4][17] = 1; doodle_sprite[0][4][18] = 1; doodle_sprite[0][4][19] = 1; doodle_sprite[0][4][20] = 1; doodle_sprite[0][4][21] = 1; doodle_sprite[0][4][22] = 1; doodle_sprite[0][4][23] = 1; doodle_sprite[0][4][24] = 1; doodle_sprite[0][4][25] = 1; doodle_sprite[0][4][26] = 1; doodle_sprite[0][4][27] = 1; doodle_sprite[0][4][28] = 1; doodle_sprite[0][4][29] = 1; doodle_sprite[0][4][30] = 1; doodle_sprite[0][4][31] = 1; doodle_sprite[0][4][32] = 1; doodle_sprite[0][4][33] = 1; doodle_sprite[0][4][34] = 1; doodle_sprite[0][4][35] = 1; doodle_sprite[0][4][36] = 1; doodle_sprite[0][4][37] = 1; doodle_sprite[0][4][38] = 1; doodle_sprite[0][4][39] = 1; doodle_sprite[0][4][40] = 1; doodle_sprite[0][4][41] = 1; doodle_sprite[0][4][42] = 1; doodle_sprite[0][4][43] = 1; doodle_sprite[0][4][44] = 1; doodle_sprite[0][4][45] = 1; doodle_sprite[0][4][46] = 1; doodle_sprite[0][4][47] = 1; doodle_sprite[0][4][48] = 1; doodle_sprite[0][4][49] = 1; doodle_sprite[0][4][50] = 1; doodle_sprite[0][4][51] = 1; doodle_sprite[0][4][52] = 1; doodle_sprite[0][4][53] = 1; doodle_sprite[0][4][54] = 1; doodle_sprite[0][4][55] = 1; doodle_sprite[0][4][56] = 1; doodle_sprite[0][4][57] = 2; doodle_sprite[0][4][58] = 2; doodle_sprite[0][4][59] = 2; doodle_sprite[0][5][16] = 2; doodle_sprite[0][5][17] = 1; doodle_sprite[0][5][18] = 1; doodle_sprite[0][5][19] = 1; doodle_sprite[0][5][20] = 1; doodle_sprite[0][5][21] = 1; doodle_sprite[0][5][22] = 1; doodle_sprite[0][5][23] = 1; doodle_sprite[0][5][24] = 1; doodle_sprite[0][5][25] = 1; doodle_sprite[0][5][26] = 1; doodle_sprite[0][5][27] = 1; doodle_sprite[0][5][28] = 1; doodle_sprite[0][5][29] = 1; doodle_sprite[0][5][30] = 1; doodle_sprite[0][5][31] = 1; doodle_sprite[0][5][32] = 1; doodle_sprite[0][5][33] = 1; doodle_sprite[0][5][34] = 1; doodle_sprite[0][5][35] = 1; doodle_sprite[0][5][36] = 1; doodle_sprite[0][5][37] = 1; doodle_sprite[0][5][38] = 1; doodle_sprite[0][5][39] = 1; doodle_sprite[0][5][40] = 1; doodle_sprite[0][5][41] = 1; doodle_sprite[0][5][42] = 1; doodle_sprite[0][5][43] = 1; doodle_sprite[0][5][44] = 1; doodle_sprite[0][5][45] = 1; doodle_sprite[0][5][46] = 1; doodle_sprite[0][5][47] = 1; doodle_sprite[0][5][48] = 1; doodle_sprite[0][5][49] = 1; doodle_sprite[0][5][50] = 1; doodle_sprite[0][5][51] = 1; doodle_sprite[0][5][52] = 1; doodle_sprite[0][5][53] = 1; doodle_sprite[0][5][54] = 1; doodle_sprite[0][5][55] = 1; doodle_sprite[0][5][56] = 1; doodle_sprite[0][5][57] = 1; doodle_sprite[0][5][58] = 1; doodle_sprite[0][5][59] = 1; doodle_sprite[0][6][16] = 2; doodle_sprite[0][6][17] = 1; doodle_sprite[0][6][18] = 1; doodle_sprite[0][6][19] = 1; doodle_sprite[0][6][20] = 1; doodle_sprite[0][6][21] = 1; doodle_sprite[0][6][22] = 1; doodle_sprite[0][6][23] = 1; doodle_sprite[0][6][24] = 1; doodle_sprite[0][6][25] = 1; doodle_sprite[0][6][26] = 1; doodle_sprite[0][6][27] = 1; doodle_sprite[0][6][28] = 1; doodle_sprite[0][6][29] = 1; doodle_sprite[0][6][30] = 1; doodle_sprite[0][6][31] = 1; doodle_sprite[0][6][32] = 1; doodle_sprite[0][6][33] = 1; doodle_sprite[0][6][34] = 1; doodle_sprite[0][6][35] = 1; doodle_sprite[0][6][36] = 1; doodle_sprite[0][6][37] = 1; doodle_sprite[0][6][38] = 1; doodle_sprite[0][6][39] = 1; doodle_sprite[0][6][40] = 1; doodle_sprite[0][6][41] = 1; doodle_sprite[0][6][42] = 1; doodle_sprite[0][6][43] = 1; doodle_sprite[0][6][44] = 1; doodle_sprite[0][6][45] = 1; doodle_sprite[0][6][46] = 1; doodle_sprite[0][6][47] = 1; doodle_sprite[0][6][48] = 1; doodle_sprite[0][6][49] = 1; doodle_sprite[0][6][50] = 1; doodle_sprite[0][6][51] = 1; doodle_sprite[0][6][52] = 1; doodle_sprite[0][6][53] = 1; doodle_sprite[0][6][54] = 1; doodle_sprite[0][6][55] = 1; doodle_sprite[0][6][56] = 1; doodle_sprite[0][6][57] = 1; doodle_sprite[0][6][58] = 1; doodle_sprite[0][6][59] = 1; doodle_sprite[0][7][16] = 2; doodle_sprite[0][7][17] = 1; doodle_sprite[0][7][18] = 1; doodle_sprite[0][7][19] = 1; doodle_sprite[0][7][20] = 1; doodle_sprite[0][7][21] = 1; doodle_sprite[0][7][22] = 1; doodle_sprite[0][7][23] = 1; doodle_sprite[0][7][24] = 1; doodle_sprite[0][7][25] = 1; doodle_sprite[0][7][26] = 1; doodle_sprite[0][7][27] = 1; doodle_sprite[0][7][28] = 1; doodle_sprite[0][7][29] = 1; doodle_sprite[0][7][30] = 1; doodle_sprite[0][7][31] = 1; doodle_sprite[0][7][32] = 1; doodle_sprite[0][7][33] = 1; doodle_sprite[0][7][34] = 1; doodle_sprite[0][7][35] = 1; doodle_sprite[0][7][36] = 1; doodle_sprite[0][7][37] = 1; doodle_sprite[0][7][38] = 1; doodle_sprite[0][7][39] = 1; doodle_sprite[0][7][40] = 1; doodle_sprite[0][7][41] = 1; doodle_sprite[0][7][42] = 1; doodle_sprite[0][7][43] = 1; doodle_sprite[0][7][44] = 1; doodle_sprite[0][7][45] = 1; doodle_sprite[0][7][46] = 1; doodle_sprite[0][7][47] = 1; doodle_sprite[0][7][48] = 1; doodle_sprite[0][7][49] = 1; doodle_sprite[0][7][50] = 1; doodle_sprite[0][7][51] = 1; doodle_sprite[0][7][52] = 1; doodle_sprite[0][7][53] = 1; doodle_sprite[0][7][54] = 1; doodle_sprite[0][7][55] = 1; doodle_sprite[0][7][56] = 1; doodle_sprite[0][7][57] = 1; doodle_sprite[0][7][58] = 1; doodle_sprite[0][7][59] = 1; doodle_sprite[0][8][12] = 2; doodle_sprite[0][8][13] = 2; doodle_sprite[0][8][14] = 2; doodle_sprite[0][8][15] = 2; doodle_sprite[0][8][16] = 2; doodle_sprite[0][8][44] = 1; doodle_sprite[0][8][45] = 1; doodle_sprite[0][8][46] = 1; doodle_sprite[0][8][47] = 1; doodle_sprite[0][8][56] = 1; doodle_sprite[0][8][57] = 1; doodle_sprite[0][8][58] = 1; doodle_sprite[0][8][59] = 1; doodle_sprite[0][8][60] = 2; doodle_sprite[0][8][61] = 1; doodle_sprite[0][8][62] = 1; doodle_sprite[0][8][63] = 1; doodle_sprite[0][8][64] = 1; doodle_sprite[0][8][65] = 2; doodle_sprite[0][8][66] = 2; doodle_sprite[0][8][67] = 2; doodle_sprite[0][8][68] = 2; doodle_sprite[0][8][69] = 2; doodle_sprite[0][8][70] = 2; doodle_sprite[0][8][71] = 2; doodle_sprite[0][9][12] = 2; doodle_sprite[0][9][13] = 2; doodle_sprite[0][9][14] = 2; doodle_sprite[0][9][15] = 2; doodle_sprite[0][9][44] = 1; doodle_sprite[0][9][45] = 1; doodle_sprite[0][9][46] = 1; doodle_sprite[0][9][47] = 1; doodle_sprite[0][9][56] = 1; doodle_sprite[0][9][57] = 1; doodle_sprite[0][9][58] = 1; doodle_sprite[0][9][59] = 1; doodle_sprite[0][9][60] = 2; doodle_sprite[0][9][61] = 1; doodle_sprite[0][9][62] = 1; doodle_sprite[0][9][63] = 1; doodle_sprite[0][9][64] = 1; doodle_sprite[0][9][65] = 2; doodle_sprite[0][9][66] = 2; doodle_sprite[0][9][67] = 2; doodle_sprite[0][9][68] = 2; doodle_sprite[0][9][69] = 2; doodle_sprite[0][9][70] = 2; doodle_sprite[0][9][71] = 2; doodle_sprite[0][10][12] = 2; doodle_sprite[0][10][13] = 2; doodle_sprite[0][10][14] = 2; doodle_sprite[0][10][15] = 2; doodle_sprite[0][10][44] = 1; doodle_sprite[0][10][45] = 1; doodle_sprite[0][10][46] = 1; doodle_sprite[0][10][47] = 1; doodle_sprite[0][10][56] = 1; doodle_sprite[0][10][57] = 1; doodle_sprite[0][10][58] = 1; doodle_sprite[0][10][59] = 1; doodle_sprite[0][10][60] = 2; doodle_sprite[0][10][61] = 1; doodle_sprite[0][10][62] = 1; doodle_sprite[0][10][63] = 1; doodle_sprite[0][10][64] = 1; doodle_sprite[0][10][65] = 2; doodle_sprite[0][10][66] = 2; doodle_sprite[0][10][67] = 2; doodle_sprite[0][10][68] = 2; doodle_sprite[0][10][69] = 2; doodle_sprite[0][10][70] = 2; doodle_sprite[0][10][71] = 2; doodle_sprite[0][11][12] = 2; doodle_sprite[0][11][13] = 2; doodle_sprite[0][11][14] = 2; doodle_sprite[0][11][15] = 1; doodle_sprite[0][11][44] = 1; doodle_sprite[0][11][45] = 1; doodle_sprite[0][11][46] = 1; doodle_sprite[0][11][47] = 1; doodle_sprite[0][11][56] = 1; doodle_sprite[0][11][57] = 1; doodle_sprite[0][11][58] = 1; doodle_sprite[0][11][59] = 1; doodle_sprite[0][11][60] = 2; doodle_sprite[0][11][61] = 1; doodle_sprite[0][11][62] = 1; doodle_sprite[0][11][63] = 1; doodle_sprite[0][11][64] = 1; doodle_sprite[0][11][65] = 2; doodle_sprite[0][11][66] = 2; doodle_sprite[0][11][67] = 2; doodle_sprite[0][11][68] = 2; doodle_sprite[0][11][69] = 2; doodle_sprite[0][11][70] = 2; doodle_sprite[0][11][71] = 2; doodle_sprite[0][12][8] = 1; doodle_sprite[0][12][9] = 1; doodle_sprite[0][12][10] = 1; doodle_sprite[0][12][11] = 1; doodle_sprite[0][12][44] = 1; doodle_sprite[0][12][45] = 1; doodle_sprite[0][12][46] = 1; doodle_sprite[0][12][47] = 1; doodle_sprite[0][12][56] = 1; doodle_sprite[0][12][57] = 1; doodle_sprite[0][12][58] = 1; doodle_sprite[0][12][59] = 1; doodle_sprite[0][12][68] = 2; doodle_sprite[0][12][69] = 2; doodle_sprite[0][12][70] = 2; doodle_sprite[0][12][71] = 2; doodle_sprite[0][13][8] = 1; doodle_sprite[0][13][9] = 1; doodle_sprite[0][13][10] = 1; doodle_sprite[0][13][11] = 1; doodle_sprite[0][13][44] = 1; doodle_sprite[0][13][45] = 1; doodle_sprite[0][13][46] = 1; doodle_sprite[0][13][47] = 1; doodle_sprite[0][13][56] = 1; doodle_sprite[0][13][57] = 1; doodle_sprite[0][13][58] = 1; doodle_sprite[0][13][59] = 1; doodle_sprite[0][13][68] = 2; doodle_sprite[0][13][69] = 2; doodle_sprite[0][13][70] = 2; doodle_sprite[0][13][71] = 2; doodle_sprite[0][14][8] = 1; doodle_sprite[0][14][9] = 1; doodle_sprite[0][14][10] = 1; doodle_sprite[0][14][11] = 1; doodle_sprite[0][14][44] = 1; doodle_sprite[0][14][45] = 1; doodle_sprite[0][14][46] = 1; doodle_sprite[0][14][47] = 1; doodle_sprite[0][14][56] = 1; doodle_sprite[0][14][57] = 1; doodle_sprite[0][14][58] = 1; doodle_sprite[0][14][59] = 1; doodle_sprite[0][14][68] = 2; doodle_sprite[0][14][69] = 2; doodle_sprite[0][14][70] = 2; doodle_sprite[0][14][71] = 2; doodle_sprite[0][15][8] = 1; doodle_sprite[0][15][9] = 1; doodle_sprite[0][15][10] = 1; doodle_sprite[0][15][11] = 1; doodle_sprite[0][15][44] = 1; doodle_sprite[0][15][45] = 1; doodle_sprite[0][15][46] = 1; doodle_sprite[0][15][47] = 1; doodle_sprite[0][15][56] = 1; doodle_sprite[0][15][57] = 1; doodle_sprite[0][15][58] = 1; doodle_sprite[0][15][59] = 1; doodle_sprite[0][15][68] = 2; doodle_sprite[0][15][69] = 2; doodle_sprite[0][15][70] = 2; doodle_sprite[0][15][71] = 2; doodle_sprite[0][16][8] = 2; doodle_sprite[0][16][9] = 2; doodle_sprite[0][16][10] = 2; doodle_sprite[0][16][11] = 1; doodle_sprite[0][16][44] = 1; doodle_sprite[0][16][45] = 1; doodle_sprite[0][16][46] = 1; doodle_sprite[0][16][47] = 1; doodle_sprite[0][16][56] = 1; doodle_sprite[0][16][57] = 1; doodle_sprite[0][16][58] = 1; doodle_sprite[0][16][59] = 1; doodle_sprite[0][17][8] = 2; doodle_sprite[0][17][9] = 2; doodle_sprite[0][17][10] = 2; doodle_sprite[0][17][11] = 1; doodle_sprite[0][17][44] = 1; doodle_sprite[0][17][45] = 1; doodle_sprite[0][17][46] = 1; doodle_sprite[0][17][47] = 1; doodle_sprite[0][17][56] = 1; doodle_sprite[0][17][57] = 1; doodle_sprite[0][17][58] = 1; doodle_sprite[0][17][59] = 1; doodle_sprite[0][18][8] = 2; doodle_sprite[0][18][9] = 2; doodle_sprite[0][18][10] = 2; doodle_sprite[0][18][11] = 1; doodle_sprite[0][18][44] = 1; doodle_sprite[0][18][45] = 1; doodle_sprite[0][18][46] = 1; doodle_sprite[0][18][47] = 1; doodle_sprite[0][18][56] = 1; doodle_sprite[0][18][57] = 1; doodle_sprite[0][18][58] = 1; doodle_sprite[0][18][59] = 1; doodle_sprite[0][19][8] = 2; doodle_sprite[0][19][9] = 2; doodle_sprite[0][19][10] = 2; doodle_sprite[0][19][11] = 1; doodle_sprite[0][19][44] = 1; doodle_sprite[0][19][45] = 1; doodle_sprite[0][19][46] = 1; doodle_sprite[0][19][47] = 1; doodle_sprite[0][19][56] = 1; doodle_sprite[0][19][57] = 1; doodle_sprite[0][19][58] = 1; doodle_sprite[0][19][59] = 1; doodle_sprite[0][20][8] = 2; doodle_sprite[0][20][9] = 2; doodle_sprite[0][20][10] = 2; doodle_sprite[0][20][11] = 1; doodle_sprite[0][20][44] = 1; doodle_sprite[0][20][45] = 1; doodle_sprite[0][20][46] = 1; doodle_sprite[0][20][47] = 1; doodle_sprite[0][20][56] = 1; doodle_sprite[0][20][57] = 1; doodle_sprite[0][20][58] = 1; doodle_sprite[0][20][59] = 1; doodle_sprite[0][20][60] = 2; doodle_sprite[0][20][61] = 2; doodle_sprite[0][20][62] = 2; doodle_sprite[0][20][63] = 1; doodle_sprite[0][20][64] = 2; doodle_sprite[0][20][65] = 2; doodle_sprite[0][20][66] = 1; doodle_sprite[0][20][67] = 2; doodle_sprite[0][20][68] = 1; doodle_sprite[0][20][69] = 1; doodle_sprite[0][20][70] = 2; doodle_sprite[0][20][71] = 2; doodle_sprite[0][21][8] = 1; doodle_sprite[0][21][9] = 1; doodle_sprite[0][21][10] = 1; doodle_sprite[0][21][11] = 1; doodle_sprite[0][21][44] = 1; doodle_sprite[0][21][45] = 1; doodle_sprite[0][21][46] = 1; doodle_sprite[0][21][47] = 1; doodle_sprite[0][21][56] = 1; doodle_sprite[0][21][57] = 1; doodle_sprite[0][21][58] = 1; doodle_sprite[0][21][59] = 1; doodle_sprite[0][21][60] = 2; doodle_sprite[0][21][61] = 2; doodle_sprite[0][21][62] = 2; doodle_sprite[0][21][63] = 1; doodle_sprite[0][21][64] = 2; doodle_sprite[0][21][65] = 2; doodle_sprite[0][21][66] = 1; doodle_sprite[0][21][67] = 2; doodle_sprite[0][21][68] = 1; doodle_sprite[0][21][69] = 1; doodle_sprite[0][21][70] = 2; doodle_sprite[0][21][71] = 2; doodle_sprite[0][22][8] = 1; doodle_sprite[0][22][9] = 1; doodle_sprite[0][22][10] = 1; doodle_sprite[0][22][11] = 1; doodle_sprite[0][22][44] = 1; doodle_sprite[0][22][45] = 1; doodle_sprite[0][22][46] = 1; doodle_sprite[0][22][47] = 1; doodle_sprite[0][22][56] = 1; doodle_sprite[0][22][57] = 1; doodle_sprite[0][22][58] = 1; doodle_sprite[0][22][59] = 1; doodle_sprite[0][22][60] = 2; doodle_sprite[0][22][61] = 2; doodle_sprite[0][22][62] = 2; doodle_sprite[0][22][63] = 1; doodle_sprite[0][22][64] = 2; doodle_sprite[0][22][65] = 2; doodle_sprite[0][22][66] = 1; doodle_sprite[0][22][67] = 2; doodle_sprite[0][22][68] = 1; doodle_sprite[0][22][69] = 1; doodle_sprite[0][22][70] = 2; doodle_sprite[0][22][71] = 2; doodle_sprite[0][23][8] = 2; doodle_sprite[0][23][9] = 2; doodle_sprite[0][23][10] = 2; doodle_sprite[0][23][11] = 1; doodle_sprite[0][23][44] = 1; doodle_sprite[0][23][45] = 1; doodle_sprite[0][23][46] = 1; doodle_sprite[0][23][47] = 1; doodle_sprite[0][23][56] = 1; doodle_sprite[0][23][57] = 1; doodle_sprite[0][23][58] = 1; doodle_sprite[0][23][59] = 1; doodle_sprite[0][23][60] = 2; doodle_sprite[0][23][61] = 2; doodle_sprite[0][23][62] = 2; doodle_sprite[0][23][63] = 1; doodle_sprite[0][23][64] = 2; doodle_sprite[0][23][65] = 2; doodle_sprite[0][23][66] = 1; doodle_sprite[0][23][67] = 2; doodle_sprite[0][23][68] = 1; doodle_sprite[0][23][69] = 1; doodle_sprite[0][23][70] = 2; doodle_sprite[0][23][71] = 2; doodle_sprite[0][24][8] = 1; doodle_sprite[0][24][9] = 1; doodle_sprite[0][24][10] = 1; doodle_sprite[0][24][11] = 1; doodle_sprite[0][24][44] = 1; doodle_sprite[0][24][45] = 1; doodle_sprite[0][24][46] = 1; doodle_sprite[0][24][47] = 1; doodle_sprite[0][24][56] = 1; doodle_sprite[0][24][57] = 1; doodle_sprite[0][24][58] = 1; doodle_sprite[0][24][59] = 1; doodle_sprite[0][24][68] = 2; doodle_sprite[0][24][69] = 2; doodle_sprite[0][24][70] = 2; doodle_sprite[0][24][71] = 2; doodle_sprite[0][25][8] = 1; doodle_sprite[0][25][9] = 1; doodle_sprite[0][25][10] = 1; doodle_sprite[0][25][11] = 1; doodle_sprite[0][25][44] = 1; doodle_sprite[0][25][45] = 1; doodle_sprite[0][25][46] = 1; doodle_sprite[0][25][47] = 1; doodle_sprite[0][25][56] = 1; doodle_sprite[0][25][57] = 1; doodle_sprite[0][25][58] = 1; doodle_sprite[0][25][59] = 1; doodle_sprite[0][25][68] = 2; doodle_sprite[0][25][69] = 2; doodle_sprite[0][25][70] = 2; doodle_sprite[0][25][71] = 2; doodle_sprite[0][26][8] = 1; doodle_sprite[0][26][9] = 1; doodle_sprite[0][26][10] = 1; doodle_sprite[0][26][11] = 1; doodle_sprite[0][26][44] = 1; doodle_sprite[0][26][45] = 1; doodle_sprite[0][26][46] = 1; doodle_sprite[0][26][47] = 1; doodle_sprite[0][26][56] = 1; doodle_sprite[0][26][57] = 1; doodle_sprite[0][26][58] = 1; doodle_sprite[0][26][59] = 1; doodle_sprite[0][26][68] = 2; doodle_sprite[0][26][69] = 2; doodle_sprite[0][26][70] = 2; doodle_sprite[0][26][71] = 2; doodle_sprite[0][27][8] = 1; doodle_sprite[0][27][9] = 1; doodle_sprite[0][27][10] = 1; doodle_sprite[0][27][11] = 1; doodle_sprite[0][27][44] = 1; doodle_sprite[0][27][45] = 1; doodle_sprite[0][27][46] = 1; doodle_sprite[0][27][47] = 1; doodle_sprite[0][27][56] = 1; doodle_sprite[0][27][57] = 1; doodle_sprite[0][27][58] = 1; doodle_sprite[0][27][59] = 1; doodle_sprite[0][27][68] = 2; doodle_sprite[0][27][69] = 2; doodle_sprite[0][27][70] = 2; doodle_sprite[0][27][71] = 2; doodle_sprite[0][28][8] = 1; doodle_sprite[0][28][9] = 1; doodle_sprite[0][28][10] = 1; doodle_sprite[0][28][11] = 1; doodle_sprite[0][28][44] = 1; doodle_sprite[0][28][45] = 1; doodle_sprite[0][28][46] = 1; doodle_sprite[0][28][47] = 1; doodle_sprite[0][28][56] = 1; doodle_sprite[0][28][57] = 1; doodle_sprite[0][28][58] = 1; doodle_sprite[0][28][59] = 1; doodle_sprite[0][29][8] = 1; doodle_sprite[0][29][9] = 1; doodle_sprite[0][29][10] = 1; doodle_sprite[0][29][11] = 1; doodle_sprite[0][29][44] = 1; doodle_sprite[0][29][45] = 1; doodle_sprite[0][29][46] = 1; doodle_sprite[0][29][47] = 1; doodle_sprite[0][29][56] = 1; doodle_sprite[0][29][57] = 1; doodle_sprite[0][29][58] = 1; doodle_sprite[0][29][59] = 1; doodle_sprite[0][30][8] = 1; doodle_sprite[0][30][9] = 1; doodle_sprite[0][30][10] = 1; doodle_sprite[0][30][11] = 1; doodle_sprite[0][30][44] = 1; doodle_sprite[0][30][45] = 1; doodle_sprite[0][30][46] = 1; doodle_sprite[0][30][47] = 1; doodle_sprite[0][30][56] = 1; doodle_sprite[0][30][57] = 1; doodle_sprite[0][30][58] = 1; doodle_sprite[0][30][59] = 1; doodle_sprite[0][31][8] = 2; doodle_sprite[0][31][9] = 2; doodle_sprite[0][31][10] = 2; doodle_sprite[0][31][11] = 1; doodle_sprite[0][31][44] = 1; doodle_sprite[0][31][45] = 1; doodle_sprite[0][31][46] = 1; doodle_sprite[0][31][47] = 1; doodle_sprite[0][31][56] = 1; doodle_sprite[0][31][57] = 1; doodle_sprite[0][31][58] = 1; doodle_sprite[0][31][59] = 1; doodle_sprite[0][32][8] = 2; doodle_sprite[0][32][9] = 2; doodle_sprite[0][32][10] = 2; doodle_sprite[0][32][11] = 1; doodle_sprite[0][32][24] = 1; doodle_sprite[0][32][25] = 1; doodle_sprite[0][32][26] = 1; doodle_sprite[0][32][27] = 1; doodle_sprite[0][32][44] = 1; doodle_sprite[0][32][45] = 1; doodle_sprite[0][32][46] = 1; doodle_sprite[0][32][47] = 1; doodle_sprite[0][32][56] = 1; doodle_sprite[0][32][57] = 1; doodle_sprite[0][32][58] = 1; doodle_sprite[0][32][59] = 1; doodle_sprite[0][32][60] = 2; doodle_sprite[0][32][61] = 2; doodle_sprite[0][32][62] = 2; doodle_sprite[0][32][63] = 2; doodle_sprite[0][32][64] = 2; doodle_sprite[0][32][65] = 2; doodle_sprite[0][32][66] = 2; doodle_sprite[0][32][67] = 2; doodle_sprite[0][32][68] = 2; doodle_sprite[0][32][69] = 2; doodle_sprite[0][32][70] = 2; doodle_sprite[0][32][71] = 2; doodle_sprite[0][33][8] = 2; doodle_sprite[0][33][9] = 2; doodle_sprite[0][33][10] = 2; doodle_sprite[0][33][11] = 1; doodle_sprite[0][33][24] = 1; doodle_sprite[0][33][25] = 1; doodle_sprite[0][33][26] = 1; doodle_sprite[0][33][27] = 1; doodle_sprite[0][33][44] = 1; doodle_sprite[0][33][45] = 1; doodle_sprite[0][33][46] = 1; doodle_sprite[0][33][47] = 1; doodle_sprite[0][33][56] = 1; doodle_sprite[0][33][57] = 1; doodle_sprite[0][33][58] = 1; doodle_sprite[0][33][59] = 1; doodle_sprite[0][33][60] = 2; doodle_sprite[0][33][61] = 2; doodle_sprite[0][33][62] = 2; doodle_sprite[0][33][63] = 2; doodle_sprite[0][33][64] = 2; doodle_sprite[0][33][65] = 2; doodle_sprite[0][33][66] = 2; doodle_sprite[0][33][67] = 2; doodle_sprite[0][33][68] = 2; doodle_sprite[0][33][69] = 2; doodle_sprite[0][33][70] = 2; doodle_sprite[0][33][71] = 2; doodle_sprite[0][34][8] = 2; doodle_sprite[0][34][9] = 2; doodle_sprite[0][34][10] = 2; doodle_sprite[0][34][11] = 1; doodle_sprite[0][34][24] = 1; doodle_sprite[0][34][25] = 1; doodle_sprite[0][34][26] = 1; doodle_sprite[0][34][27] = 1; doodle_sprite[0][34][44] = 1; doodle_sprite[0][34][45] = 1; doodle_sprite[0][34][46] = 1; doodle_sprite[0][34][47] = 1; doodle_sprite[0][34][56] = 1; doodle_sprite[0][34][57] = 1; doodle_sprite[0][34][58] = 1; doodle_sprite[0][34][59] = 1; doodle_sprite[0][34][60] = 2; doodle_sprite[0][34][61] = 2; doodle_sprite[0][34][62] = 2; doodle_sprite[0][34][63] = 2; doodle_sprite[0][34][64] = 2; doodle_sprite[0][34][65] = 2; doodle_sprite[0][34][66] = 2; doodle_sprite[0][34][67] = 2; doodle_sprite[0][34][68] = 2; doodle_sprite[0][34][69] = 2; doodle_sprite[0][34][70] = 2; doodle_sprite[0][34][71] = 2; doodle_sprite[0][35][8] = 2; doodle_sprite[0][35][9] = 2; doodle_sprite[0][35][10] = 2; doodle_sprite[0][35][11] = 1; doodle_sprite[0][35][24] = 1; doodle_sprite[0][35][25] = 1; doodle_sprite[0][35][26] = 1; doodle_sprite[0][35][27] = 1; doodle_sprite[0][35][44] = 1; doodle_sprite[0][35][45] = 1; doodle_sprite[0][35][46] = 1; doodle_sprite[0][35][47] = 1; doodle_sprite[0][35][56] = 1; doodle_sprite[0][35][57] = 1; doodle_sprite[0][35][58] = 1; doodle_sprite[0][35][59] = 1; doodle_sprite[0][35][60] = 2; doodle_sprite[0][35][61] = 2; doodle_sprite[0][35][62] = 2; doodle_sprite[0][35][63] = 2; doodle_sprite[0][35][64] = 2; doodle_sprite[0][35][65] = 2; doodle_sprite[0][35][66] = 2; doodle_sprite[0][35][67] = 2; doodle_sprite[0][35][68] = 2; doodle_sprite[0][35][69] = 2; doodle_sprite[0][35][70] = 2; doodle_sprite[0][35][71] = 2; doodle_sprite[0][36][8] = 2; doodle_sprite[0][36][9] = 2; doodle_sprite[0][36][10] = 2; doodle_sprite[0][36][11] = 1; doodle_sprite[0][36][44] = 1; doodle_sprite[0][36][45] = 1; doodle_sprite[0][36][46] = 1; doodle_sprite[0][36][47] = 1; doodle_sprite[0][36][56] = 1; doodle_sprite[0][36][57] = 1; doodle_sprite[0][36][58] = 1; doodle_sprite[0][36][59] = 1; doodle_sprite[0][36][68] = 2; doodle_sprite[0][36][69] = 2; doodle_sprite[0][36][70] = 2; doodle_sprite[0][36][71] = 2; doodle_sprite[0][37][8] = 2; doodle_sprite[0][37][9] = 2; doodle_sprite[0][37][10] = 2; doodle_sprite[0][37][11] = 1; doodle_sprite[0][37][44] = 1; doodle_sprite[0][37][45] = 1; doodle_sprite[0][37][46] = 1; doodle_sprite[0][37][47] = 1; doodle_sprite[0][37][56] = 1; doodle_sprite[0][37][57] = 1; doodle_sprite[0][37][58] = 1; doodle_sprite[0][37][59] = 1; doodle_sprite[0][37][68] = 2; doodle_sprite[0][37][69] = 2; doodle_sprite[0][37][70] = 2; doodle_sprite[0][37][71] = 2; doodle_sprite[0][38][8] = 2; doodle_sprite[0][38][9] = 2; doodle_sprite[0][38][10] = 2; doodle_sprite[0][38][11] = 2; doodle_sprite[0][38][44] = 1; doodle_sprite[0][38][45] = 1; doodle_sprite[0][38][46] = 1; doodle_sprite[0][38][47] = 1; doodle_sprite[0][38][56] = 1; doodle_sprite[0][38][57] = 1; doodle_sprite[0][38][58] = 1; doodle_sprite[0][38][59] = 1; doodle_sprite[0][38][68] = 2; doodle_sprite[0][38][69] = 2; doodle_sprite[0][38][70] = 2; doodle_sprite[0][38][71] = 2; doodle_sprite[0][39][8] = 2; doodle_sprite[0][39][9] = 2; doodle_sprite[0][39][10] = 2; doodle_sprite[0][39][11] = 2; doodle_sprite[0][39][44] = 1; doodle_sprite[0][39][45] = 1; doodle_sprite[0][39][46] = 1; doodle_sprite[0][39][47] = 1; doodle_sprite[0][39][56] = 1; doodle_sprite[0][39][57] = 1; doodle_sprite[0][39][58] = 1; doodle_sprite[0][39][59] = 1; doodle_sprite[0][39][68] = 2; doodle_sprite[0][39][69] = 2; doodle_sprite[0][39][70] = 2; doodle_sprite[0][39][71] = 2; doodle_sprite[0][40][8] = 2; doodle_sprite[0][40][9] = 2; doodle_sprite[0][40][10] = 2; doodle_sprite[0][40][11] = 2; doodle_sprite[0][40][24] = 1; doodle_sprite[0][40][25] = 1; doodle_sprite[0][40][26] = 1; doodle_sprite[0][40][27] = 1; doodle_sprite[0][40][44] = 1; doodle_sprite[0][40][45] = 1; doodle_sprite[0][40][46] = 1; doodle_sprite[0][40][47] = 1; doodle_sprite[0][40][56] = 1; doodle_sprite[0][40][57] = 1; doodle_sprite[0][40][58] = 1; doodle_sprite[0][40][59] = 1; doodle_sprite[0][41][8] = 2; doodle_sprite[0][41][9] = 2; doodle_sprite[0][41][10] = 2; doodle_sprite[0][41][11] = 2; doodle_sprite[0][41][24] = 1; doodle_sprite[0][41][25] = 1; doodle_sprite[0][41][26] = 1; doodle_sprite[0][41][27] = 1; doodle_sprite[0][41][44] = 1; doodle_sprite[0][41][45] = 1; doodle_sprite[0][41][46] = 1; doodle_sprite[0][41][47] = 1; doodle_sprite[0][41][56] = 1; doodle_sprite[0][41][57] = 1; doodle_sprite[0][41][58] = 1; doodle_sprite[0][41][59] = 1; doodle_sprite[0][42][8] = 2; doodle_sprite[0][42][9] = 2; doodle_sprite[0][42][10] = 2; doodle_sprite[0][42][11] = 2; doodle_sprite[0][42][24] = 1; doodle_sprite[0][42][25] = 1; doodle_sprite[0][42][26] = 1; doodle_sprite[0][42][27] = 1; doodle_sprite[0][42][44] = 1; doodle_sprite[0][42][45] = 1; doodle_sprite[0][42][46] = 1; doodle_sprite[0][42][47] = 1; doodle_sprite[0][42][56] = 1; doodle_sprite[0][42][57] = 1; doodle_sprite[0][42][58] = 1; doodle_sprite[0][42][59] = 1; doodle_sprite[0][43][8] = 2; doodle_sprite[0][43][9] = 2; doodle_sprite[0][43][10] = 2; doodle_sprite[0][43][11] = 2; doodle_sprite[0][43][24] = 1; doodle_sprite[0][43][25] = 1; doodle_sprite[0][43][26] = 1; doodle_sprite[0][43][27] = 1; doodle_sprite[0][43][44] = 1; doodle_sprite[0][43][45] = 1; doodle_sprite[0][43][46] = 1; doodle_sprite[0][43][47] = 1; doodle_sprite[0][43][56] = 1; doodle_sprite[0][43][57] = 1; doodle_sprite[0][43][58] = 1; doodle_sprite[0][43][59] = 1; doodle_sprite[0][44][12] = 2; doodle_sprite[0][44][13] = 2; doodle_sprite[0][44][14] = 2; doodle_sprite[0][44][15] = 2; doodle_sprite[0][44][16] = 2; doodle_sprite[0][44][44] = 1; doodle_sprite[0][44][45] = 1; doodle_sprite[0][44][46] = 1; doodle_sprite[0][44][47] = 1; doodle_sprite[0][44][56] = 1; doodle_sprite[0][44][57] = 1; doodle_sprite[0][44][58] = 1; doodle_sprite[0][44][59] = 1; doodle_sprite[0][44][60] = 2; doodle_sprite[0][44][61] = 2; doodle_sprite[0][44][62] = 2; doodle_sprite[0][44][63] = 2; doodle_sprite[0][44][64] = 2; doodle_sprite[0][44][65] = 2; doodle_sprite[0][44][66] = 2; doodle_sprite[0][44][67] = 2; doodle_sprite[0][44][68] = 2; doodle_sprite[0][44][69] = 2; doodle_sprite[0][44][70] = 2; doodle_sprite[0][44][71] = 2; doodle_sprite[0][45][12] = 2; doodle_sprite[0][45][13] = 2; doodle_sprite[0][45][14] = 2; doodle_sprite[0][45][15] = 2; doodle_sprite[0][45][16] = 2; doodle_sprite[0][45][44] = 1; doodle_sprite[0][45][45] = 1; doodle_sprite[0][45][46] = 1; doodle_sprite[0][45][47] = 1; doodle_sprite[0][45][56] = 1; doodle_sprite[0][45][57] = 1; doodle_sprite[0][45][58] = 1; doodle_sprite[0][45][59] = 1; doodle_sprite[0][45][60] = 2; doodle_sprite[0][45][61] = 2; doodle_sprite[0][45][62] = 2; doodle_sprite[0][45][63] = 2; doodle_sprite[0][45][64] = 2; doodle_sprite[0][45][65] = 2; doodle_sprite[0][45][66] = 2; doodle_sprite[0][45][67] = 2; doodle_sprite[0][45][68] = 2; doodle_sprite[0][45][69] = 2; doodle_sprite[0][45][70] = 2; doodle_sprite[0][45][71] = 2; doodle_sprite[0][46][12] = 2; doodle_sprite[0][46][13] = 2; doodle_sprite[0][46][14] = 2; doodle_sprite[0][46][15] = 2; doodle_sprite[0][46][16] = 2; doodle_sprite[0][46][44] = 1; doodle_sprite[0][46][45] = 1; doodle_sprite[0][46][46] = 1; doodle_sprite[0][46][47] = 1; doodle_sprite[0][46][56] = 1; doodle_sprite[0][46][57] = 1; doodle_sprite[0][46][58] = 1; doodle_sprite[0][46][59] = 1; doodle_sprite[0][46][60] = 2; doodle_sprite[0][46][61] = 2; doodle_sprite[0][46][62] = 2; doodle_sprite[0][46][63] = 2; doodle_sprite[0][46][64] = 2; doodle_sprite[0][46][65] = 2; doodle_sprite[0][46][66] = 2; doodle_sprite[0][46][67] = 2; doodle_sprite[0][46][68] = 2; doodle_sprite[0][46][69] = 2; doodle_sprite[0][46][70] = 2; doodle_sprite[0][46][71] = 2; doodle_sprite[0][47][12] = 2; doodle_sprite[0][47][13] = 2; doodle_sprite[0][47][14] = 2; doodle_sprite[0][47][15] = 2; doodle_sprite[0][47][16] = 2; doodle_sprite[0][47][44] = 1; doodle_sprite[0][47][45] = 1; doodle_sprite[0][47][46] = 1; doodle_sprite[0][47][47] = 1; doodle_sprite[0][47][56] = 1; doodle_sprite[0][47][57] = 1; doodle_sprite[0][47][58] = 1; doodle_sprite[0][47][59] = 1; doodle_sprite[0][47][60] = 2; doodle_sprite[0][47][61] = 2; doodle_sprite[0][47][62] = 2; doodle_sprite[0][47][63] = 2; doodle_sprite[0][47][64] = 2; doodle_sprite[0][47][65] = 2; doodle_sprite[0][47][66] = 2; doodle_sprite[0][47][67] = 2; doodle_sprite[0][47][68] = 2; doodle_sprite[0][47][69] = 2; doodle_sprite[0][47][70] = 2; doodle_sprite[0][47][71] = 2; doodle_sprite[0][48][16] = 2; doodle_sprite[0][48][17] = 2; doodle_sprite[0][48][18] = 2; doodle_sprite[0][48][19] = 2; doodle_sprite[0][48][20] = 2; doodle_sprite[0][48][21] = 2; doodle_sprite[0][48][22] = 2; doodle_sprite[0][48][23] = 2; doodle_sprite[0][48][24] = 2; doodle_sprite[0][48][25] = 2; doodle_sprite[0][48][26] = 2; doodle_sprite[0][48][27] = 1; doodle_sprite[0][48][36] = 1; doodle_sprite[0][48][37] = 1; doodle_sprite[0][48][38] = 1; doodle_sprite[0][48][39] = 1; doodle_sprite[0][48][40] = 1; doodle_sprite[0][48][41] = 1; doodle_sprite[0][48][42] = 1; doodle_sprite[0][48][43] = 1; doodle_sprite[0][48][44] = 1; doodle_sprite[0][48][45] = 1; doodle_sprite[0][48][46] = 1; doodle_sprite[0][48][47] = 1; doodle_sprite[0][48][48] = 1; doodle_sprite[0][48][49] = 1; doodle_sprite[0][48][50] = 1; doodle_sprite[0][48][51] = 1; doodle_sprite[0][48][52] = 1; doodle_sprite[0][48][53] = 1; doodle_sprite[0][48][54] = 1; doodle_sprite[0][48][55] = 1; doodle_sprite[0][48][56] = 1; doodle_sprite[0][48][57] = 1; doodle_sprite[0][48][58] = 1; doodle_sprite[0][48][59] = 1; doodle_sprite[0][48][68] = 2; doodle_sprite[0][48][69] = 2; doodle_sprite[0][48][70] = 2; doodle_sprite[0][48][71] = 2; doodle_sprite[0][49][16] = 2; doodle_sprite[0][49][17] = 2; doodle_sprite[0][49][18] = 2; doodle_sprite[0][49][19] = 2; doodle_sprite[0][49][20] = 2; doodle_sprite[0][49][21] = 2; doodle_sprite[0][49][22] = 2; doodle_sprite[0][49][23] = 2; doodle_sprite[0][49][24] = 1; doodle_sprite[0][49][25] = 1; doodle_sprite[0][49][26] = 1; doodle_sprite[0][49][27] = 1; doodle_sprite[0][49][36] = 1; doodle_sprite[0][49][37] = 1; doodle_sprite[0][49][38] = 1; doodle_sprite[0][49][39] = 1; doodle_sprite[0][49][40] = 1; doodle_sprite[0][49][41] = 1; doodle_sprite[0][49][42] = 1; doodle_sprite[0][49][43] = 1; doodle_sprite[0][49][44] = 1; doodle_sprite[0][49][45] = 1; doodle_sprite[0][49][46] = 1; doodle_sprite[0][49][47] = 1; doodle_sprite[0][49][48] = 1; doodle_sprite[0][49][49] = 1; doodle_sprite[0][49][50] = 1; doodle_sprite[0][49][51] = 1; doodle_sprite[0][49][52] = 1; doodle_sprite[0][49][53] = 1; doodle_sprite[0][49][54] = 1; doodle_sprite[0][49][55] = 1; doodle_sprite[0][49][56] = 1; doodle_sprite[0][49][57] = 1; doodle_sprite[0][49][58] = 1; doodle_sprite[0][49][59] = 1; doodle_sprite[0][49][68] = 2; doodle_sprite[0][49][69] = 2; doodle_sprite[0][49][70] = 2; doodle_sprite[0][49][71] = 2; doodle_sprite[0][50][16] = 2; doodle_sprite[0][50][17] = 2; doodle_sprite[0][50][18] = 2; doodle_sprite[0][50][19] = 2; doodle_sprite[0][50][20] = 2; doodle_sprite[0][50][21] = 2; doodle_sprite[0][50][22] = 2; doodle_sprite[0][50][23] = 2; doodle_sprite[0][50][24] = 1; doodle_sprite[0][50][25] = 1; doodle_sprite[0][50][26] = 1; doodle_sprite[0][50][27] = 1; doodle_sprite[0][50][36] = 1; doodle_sprite[0][50][37] = 1; doodle_sprite[0][50][38] = 1; doodle_sprite[0][50][39] = 1; doodle_sprite[0][50][40] = 1; doodle_sprite[0][50][41] = 1; doodle_sprite[0][50][42] = 1; doodle_sprite[0][50][43] = 1; doodle_sprite[0][50][44] = 1; doodle_sprite[0][50][45] = 1; doodle_sprite[0][50][46] = 1; doodle_sprite[0][50][47] = 1; doodle_sprite[0][50][48] = 1; doodle_sprite[0][50][49] = 1; doodle_sprite[0][50][50] = 1; doodle_sprite[0][50][51] = 1; doodle_sprite[0][50][52] = 1; doodle_sprite[0][50][53] = 1; doodle_sprite[0][50][54] = 1; doodle_sprite[0][50][55] = 1; doodle_sprite[0][50][56] = 1; doodle_sprite[0][50][57] = 2; doodle_sprite[0][50][58] = 2; doodle_sprite[0][50][59] = 2; doodle_sprite[0][50][68] = 2; doodle_sprite[0][50][69] = 2; doodle_sprite[0][50][70] = 2; doodle_sprite[0][50][71] = 2; doodle_sprite[0][51][16] = 2; doodle_sprite[0][51][17] = 2; doodle_sprite[0][51][18] = 2; doodle_sprite[0][51][19] = 2; doodle_sprite[0][51][20] = 2; doodle_sprite[0][51][21] = 2; doodle_sprite[0][51][22] = 2; doodle_sprite[0][51][23] = 2; doodle_sprite[0][51][24] = 1; doodle_sprite[0][51][25] = 1; doodle_sprite[0][51][26] = 1; doodle_sprite[0][51][27] = 1; doodle_sprite[0][51][35] = 2; doodle_sprite[0][51][36] = 1; doodle_sprite[0][51][37] = 1; doodle_sprite[0][51][38] = 1; doodle_sprite[0][51][39] = 1; doodle_sprite[0][51][40] = 1; doodle_sprite[0][51][41] = 1; doodle_sprite[0][51][42] = 1; doodle_sprite[0][51][43] = 1; doodle_sprite[0][51][44] = 1; doodle_sprite[0][51][45] = 1; doodle_sprite[0][51][46] = 1; doodle_sprite[0][51][47] = 1; doodle_sprite[0][51][48] = 1; doodle_sprite[0][51][49] = 1; doodle_sprite[0][51][50] = 1; doodle_sprite[0][51][51] = 1; doodle_sprite[0][51][52] = 1; doodle_sprite[0][51][53] = 1; doodle_sprite[0][51][54] = 1; doodle_sprite[0][51][55] = 1; doodle_sprite[0][51][56] = 1; doodle_sprite[0][51][57] = 2; doodle_sprite[0][51][58] = 2; doodle_sprite[0][51][59] = 2; doodle_sprite[0][51][68] = 2; doodle_sprite[0][51][69] = 2; doodle_sprite[0][51][70] = 2; doodle_sprite[0][51][71] = 2; doodle_sprite[0][52][24] = 1; doodle_sprite[0][52][25] = 1; doodle_sprite[0][52][26] = 1; doodle_sprite[0][52][27] = 1; doodle_sprite[0][52][32] = 1; doodle_sprite[0][52][33] = 1; doodle_sprite[0][52][34] = 1; doodle_sprite[0][52][35] = 1; doodle_sprite[0][53][24] = 1; doodle_sprite[0][53][25] = 1; doodle_sprite[0][53][26] = 1; doodle_sprite[0][53][27] = 1; doodle_sprite[0][53][32] = 1; doodle_sprite[0][53][33] = 1; doodle_sprite[0][53][34] = 1; doodle_sprite[0][53][35] = 1; doodle_sprite[0][54][24] = 1; doodle_sprite[0][54][25] = 1; doodle_sprite[0][54][26] = 1; doodle_sprite[0][54][27] = 1; doodle_sprite[0][54][32] = 1; doodle_sprite[0][54][33] = 1; doodle_sprite[0][54][34] = 1; doodle_sprite[0][54][35] = 1; doodle_sprite[0][55][24] = 1; doodle_sprite[0][55][25] = 1; doodle_sprite[0][55][26] = 1; doodle_sprite[0][55][27] = 1; doodle_sprite[0][55][32] = 1; doodle_sprite[0][55][33] = 1; doodle_sprite[0][55][34] = 1; doodle_sprite[0][55][35] = 1; doodle_sprite[0][56][24] = 1; doodle_sprite[0][56][25] = 1; doodle_sprite[0][56][26] = 1; doodle_sprite[0][56][27] = 1; doodle_sprite[0][56][32] = 1; doodle_sprite[0][56][33] = 1; doodle_sprite[0][56][34] = 1; doodle_sprite[0][56][35] = 1; doodle_sprite[0][57][24] = 1; doodle_sprite[0][57][25] = 1; doodle_sprite[0][57][26] = 1; doodle_sprite[0][57][27] = 1; doodle_sprite[0][57][32] = 1; doodle_sprite[0][57][33] = 1; doodle_sprite[0][57][34] = 1; doodle_sprite[0][57][35] = 1; doodle_sprite[0][58][24] = 1; doodle_sprite[0][58][25] = 1; doodle_sprite[0][58][26] = 1; doodle_sprite[0][58][27] = 1; doodle_sprite[0][58][32] = 1; doodle_sprite[0][58][33] = 1; doodle_sprite[0][58][34] = 1; doodle_sprite[0][58][35] = 1; doodle_sprite[0][59][24] = 1; doodle_sprite[0][59][25] = 1; doodle_sprite[0][59][26] = 1; doodle_sprite[0][59][27] = 1; doodle_sprite[0][59][32] = 1; doodle_sprite[0][59][33] = 1; doodle_sprite[0][59][34] = 1; doodle_sprite[0][59][35] = 1; doodle_sprite[0][60][24] = 1; doodle_sprite[0][60][25] = 1; doodle_sprite[0][60][26] = 1; doodle_sprite[0][60][27] = 1; doodle_sprite[0][60][32] = 1; doodle_sprite[0][60][33] = 1; doodle_sprite[0][60][34] = 1; doodle_sprite[0][60][35] = 1; doodle_sprite[0][61][24] = 1; doodle_sprite[0][61][25] = 1; doodle_sprite[0][61][26] = 1; doodle_sprite[0][61][27] = 1; doodle_sprite[0][61][32] = 1; doodle_sprite[0][61][33] = 1; doodle_sprite[0][61][34] = 1; doodle_sprite[0][61][35] = 1; doodle_sprite[0][62][24] = 1; doodle_sprite[0][62][25] = 1; doodle_sprite[0][62][26] = 1; doodle_sprite[0][62][27] = 1; doodle_sprite[0][62][32] = 1; doodle_sprite[0][62][33] = 1; doodle_sprite[0][62][34] = 1; doodle_sprite[0][62][35] = 1; doodle_sprite[0][63][24] = 1; doodle_sprite[0][63][25] = 1; doodle_sprite[0][63][26] = 1; doodle_sprite[0][63][27] = 1; doodle_sprite[0][63][32] = 1; doodle_sprite[0][63][33] = 1; doodle_sprite[0][63][34] = 1; doodle_sprite[0][63][35] = 1; doodle_sprite[0][64][24] = 1; doodle_sprite[0][64][25] = 1; doodle_sprite[0][64][26] = 1; doodle_sprite[0][64][27] = 1; doodle_sprite[0][64][28] = 1; doodle_sprite[0][64][29] = 1; doodle_sprite[0][64][30] = 1; doodle_sprite[0][64][31] = 1; doodle_sprite[0][64][32] = 1; doodle_sprite[0][64][33] = 1; doodle_sprite[0][64][34] = 1; doodle_sprite[0][64][35] = 1; doodle_sprite[0][65][24] = 1; doodle_sprite[0][65][25] = 1; doodle_sprite[0][65][26] = 1; doodle_sprite[0][65][27] = 1; doodle_sprite[0][65][28] = 1; doodle_sprite[0][65][29] = 1; doodle_sprite[0][65][30] = 1; doodle_sprite[0][65][31] = 1; doodle_sprite[0][65][32] = 1; doodle_sprite[0][65][33] = 1; doodle_sprite[0][65][34] = 1; doodle_sprite[0][65][35] = 1; doodle_sprite[0][66][24] = 1; doodle_sprite[0][66][25] = 1; doodle_sprite[0][66][26] = 1; doodle_sprite[0][66][27] = 1; doodle_sprite[0][66][28] = 1; doodle_sprite[0][66][29] = 1; doodle_sprite[0][66][30] = 1; doodle_sprite[0][66][31] = 1; doodle_sprite[0][66][32] = 1; doodle_sprite[0][66][33] = 1; doodle_sprite[0][66][34] = 1; doodle_sprite[0][66][35] = 1; doodle_sprite[0][67][24] = 1; doodle_sprite[0][67][25] = 1; doodle_sprite[0][67][26] = 1; doodle_sprite[0][67][27] = 1; doodle_sprite[0][67][28] = 1; doodle_sprite[0][67][29] = 1; doodle_sprite[0][67][30] = 1; doodle_sprite[0][67][31] = 1; doodle_sprite[0][67][32] = 1; doodle_sprite[0][67][33] = 1; doodle_sprite[0][67][34] = 1; doodle_sprite[0][67][35] = 1; doodle_sprite[0][68][24] = 2; doodle_sprite[0][68][25] = 2; doodle_sprite[0][68][26] = 2; doodle_sprite[0][68][27] = 1; doodle_sprite[0][68][32] = 1; doodle_sprite[0][68][33] = 1; doodle_sprite[0][68][34] = 1; doodle_sprite[0][68][35] = 1; doodle_sprite[0][69][24] = 2; doodle_sprite[0][69][25] = 2; doodle_sprite[0][69][26] = 2; doodle_sprite[0][69][27] = 1; doodle_sprite[0][69][32] = 1; doodle_sprite[0][69][33] = 1; doodle_sprite[0][69][34] = 1; doodle_sprite[0][69][35] = 1; doodle_sprite[0][70][24] = 2; doodle_sprite[0][70][25] = 2; doodle_sprite[0][70][26] = 2; doodle_sprite[0][70][27] = 1; doodle_sprite[0][70][32] = 1; doodle_sprite[0][70][33] = 1; doodle_sprite[0][70][34] = 1; doodle_sprite[0][70][35] = 1; doodle_sprite[0][71][24] = 2; doodle_sprite[0][71][25] = 2; doodle_sprite[0][71][26] = 2; doodle_sprite[0][71][27] = 1; doodle_sprite[0][71][32] = 1; doodle_sprite[0][71][33] = 1; doodle_sprite[0][71][34] = 1; doodle_sprite[0][71][35] = 1; doodle_sprite[0][72][24] = 2; doodle_sprite[0][72][25] = 2; doodle_sprite[0][72][26] = 2; doodle_sprite[0][72][27] = 1; doodle_sprite[0][72][28] = 1; doodle_sprite[0][72][29] = 1; doodle_sprite[0][72][30] = 1; doodle_sprite[0][72][31] = 1; doodle_sprite[0][72][32] = 1; doodle_sprite[0][72][33] = 2; doodle_sprite[0][72][34] = 2; doodle_sprite[0][72][35] = 2; doodle_sprite[0][73][24] = 2; doodle_sprite[0][73][25] = 2; doodle_sprite[0][73][26] = 2; doodle_sprite[0][73][27] = 2; doodle_sprite[0][73][28] = 2; doodle_sprite[0][73][29] = 2; doodle_sprite[0][73][30] = 2; doodle_sprite[0][73][31] = 2; doodle_sprite[0][73][32] = 2; doodle_sprite[0][73][33] = 2; doodle_sprite[0][73][34] = 2; doodle_sprite[0][73][35] = 2; doodle_sprite[0][74][24] = 2; doodle_sprite[0][74][25] = 2; doodle_sprite[0][74][26] = 2; doodle_sprite[0][74][27] = 2; doodle_sprite[0][74][28] = 2; doodle_sprite[0][74][29] = 2; doodle_sprite[0][74][30] = 2; doodle_sprite[0][74][31] = 2; doodle_sprite[0][74][32] = 2; doodle_sprite[0][74][33] = 2; doodle_sprite[0][74][34] = 2; doodle_sprite[0][74][35] = 2; doodle_sprite[0][75][24] = 2; doodle_sprite[0][75][25] = 2; doodle_sprite[0][75][26] = 2; doodle_sprite[0][75][27] = 2; doodle_sprite[0][75][28] = 2; doodle_sprite[0][75][29] = 2; doodle_sprite[0][75][30] = 2; doodle_sprite[0][75][31] = 2; doodle_sprite[0][75][32] = 2; doodle_sprite[0][75][33] = 2; doodle_sprite[0][75][34] = 2; doodle_sprite[0][75][35] = 2; 
					doodle_sprite[1][4][16] = 2; doodle_sprite[1][4][17] = 1; doodle_sprite[1][4][18] = 1; doodle_sprite[1][4][19] = 1; doodle_sprite[1][4][20] = 1; doodle_sprite[1][4][21] = 1; doodle_sprite[1][4][22] = 1; doodle_sprite[1][4][23] = 1; doodle_sprite[1][4][24] = 1; doodle_sprite[1][4][25] = 1; doodle_sprite[1][4][26] = 1; doodle_sprite[1][4][27] = 1; doodle_sprite[1][4][28] = 1; doodle_sprite[1][4][29] = 1; doodle_sprite[1][4][30] = 1; doodle_sprite[1][4][31] = 1; doodle_sprite[1][4][32] = 1; doodle_sprite[1][4][33] = 1; doodle_sprite[1][4][34] = 1; doodle_sprite[1][4][35] = 1; doodle_sprite[1][4][36] = 1; doodle_sprite[1][4][37] = 1; doodle_sprite[1][4][38] = 1; doodle_sprite[1][4][39] = 1; doodle_sprite[1][4][40] = 1; doodle_sprite[1][4][41] = 1; doodle_sprite[1][4][42] = 1; doodle_sprite[1][4][43] = 1; doodle_sprite[1][4][44] = 1; doodle_sprite[1][4][45] = 1; doodle_sprite[1][4][46] = 1; doodle_sprite[1][4][47] = 1; doodle_sprite[1][4][48] = 1; doodle_sprite[1][4][49] = 1; doodle_sprite[1][4][50] = 1; doodle_sprite[1][4][51] = 1; doodle_sprite[1][4][52] = 1; doodle_sprite[1][4][53] = 1; doodle_sprite[1][4][54] = 1; doodle_sprite[1][4][55] = 1; doodle_sprite[1][4][56] = 1; doodle_sprite[1][4][57] = 2; doodle_sprite[1][4][58] = 2; doodle_sprite[1][4][59] = 2; doodle_sprite[1][5][16] = 2; doodle_sprite[1][5][17] = 1; doodle_sprite[1][5][18] = 1; doodle_sprite[1][5][19] = 1; doodle_sprite[1][5][20] = 1; doodle_sprite[1][5][21] = 1; doodle_sprite[1][5][22] = 1; doodle_sprite[1][5][23] = 1; doodle_sprite[1][5][24] = 1; doodle_sprite[1][5][25] = 1; doodle_sprite[1][5][26] = 1; doodle_sprite[1][5][27] = 1; doodle_sprite[1][5][28] = 1; doodle_sprite[1][5][29] = 1; doodle_sprite[1][5][30] = 1; doodle_sprite[1][5][31] = 1; doodle_sprite[1][5][32] = 1; doodle_sprite[1][5][33] = 1; doodle_sprite[1][5][34] = 1; doodle_sprite[1][5][35] = 1; doodle_sprite[1][5][36] = 1; doodle_sprite[1][5][37] = 1; doodle_sprite[1][5][38] = 1; doodle_sprite[1][5][39] = 1; doodle_sprite[1][5][40] = 1; doodle_sprite[1][5][41] = 1; doodle_sprite[1][5][42] = 1; doodle_sprite[1][5][43] = 1; doodle_sprite[1][5][44] = 1; doodle_sprite[1][5][45] = 1; doodle_sprite[1][5][46] = 1; doodle_sprite[1][5][47] = 1; doodle_sprite[1][5][48] = 1; doodle_sprite[1][5][49] = 1; doodle_sprite[1][5][50] = 1; doodle_sprite[1][5][51] = 1; doodle_sprite[1][5][52] = 1; doodle_sprite[1][5][53] = 1; doodle_sprite[1][5][54] = 1; doodle_sprite[1][5][55] = 1; doodle_sprite[1][5][56] = 1; doodle_sprite[1][5][57] = 1; doodle_sprite[1][5][58] = 1; doodle_sprite[1][5][59] = 1; doodle_sprite[1][6][16] = 2; doodle_sprite[1][6][17] = 1; doodle_sprite[1][6][18] = 1; doodle_sprite[1][6][19] = 1; doodle_sprite[1][6][20] = 1; doodle_sprite[1][6][21] = 1; doodle_sprite[1][6][22] = 1; doodle_sprite[1][6][23] = 1; doodle_sprite[1][6][24] = 1; doodle_sprite[1][6][25] = 1; doodle_sprite[1][6][26] = 1; doodle_sprite[1][6][27] = 1; doodle_sprite[1][6][28] = 1; doodle_sprite[1][6][29] = 1; doodle_sprite[1][6][30] = 1; doodle_sprite[1][6][31] = 1; doodle_sprite[1][6][32] = 1; doodle_sprite[1][6][33] = 1; doodle_sprite[1][6][34] = 1; doodle_sprite[1][6][35] = 1; doodle_sprite[1][6][36] = 1; doodle_sprite[1][6][37] = 1; doodle_sprite[1][6][38] = 1; doodle_sprite[1][6][39] = 1; doodle_sprite[1][6][40] = 1; doodle_sprite[1][6][41] = 1; doodle_sprite[1][6][42] = 1; doodle_sprite[1][6][43] = 1; doodle_sprite[1][6][44] = 1; doodle_sprite[1][6][45] = 1; doodle_sprite[1][6][46] = 1; doodle_sprite[1][6][47] = 1; doodle_sprite[1][6][48] = 1; doodle_sprite[1][6][49] = 1; doodle_sprite[1][6][50] = 1; doodle_sprite[1][6][51] = 1; doodle_sprite[1][6][52] = 1; doodle_sprite[1][6][53] = 1; doodle_sprite[1][6][54] = 1; doodle_sprite[1][6][55] = 1; doodle_sprite[1][6][56] = 1; doodle_sprite[1][6][57] = 1; doodle_sprite[1][6][58] = 1; doodle_sprite[1][6][59] = 1; doodle_sprite[1][7][16] = 2; doodle_sprite[1][7][17] = 1; doodle_sprite[1][7][18] = 1; doodle_sprite[1][7][19] = 1; doodle_sprite[1][7][20] = 1; doodle_sprite[1][7][21] = 1; doodle_sprite[1][7][22] = 1; doodle_sprite[1][7][23] = 1; doodle_sprite[1][7][24] = 1; doodle_sprite[1][7][25] = 1; doodle_sprite[1][7][26] = 1; doodle_sprite[1][7][27] = 1; doodle_sprite[1][7][28] = 1; doodle_sprite[1][7][29] = 1; doodle_sprite[1][7][30] = 1; doodle_sprite[1][7][31] = 1; doodle_sprite[1][7][32] = 1; doodle_sprite[1][7][33] = 1; doodle_sprite[1][7][34] = 1; doodle_sprite[1][7][35] = 1; doodle_sprite[1][7][36] = 1; doodle_sprite[1][7][37] = 1; doodle_sprite[1][7][38] = 1; doodle_sprite[1][7][39] = 1; doodle_sprite[1][7][40] = 1; doodle_sprite[1][7][41] = 1; doodle_sprite[1][7][42] = 1; doodle_sprite[1][7][43] = 1; doodle_sprite[1][7][44] = 1; doodle_sprite[1][7][45] = 1; doodle_sprite[1][7][46] = 1; doodle_sprite[1][7][47] = 1; doodle_sprite[1][7][48] = 1; doodle_sprite[1][7][49] = 1; doodle_sprite[1][7][50] = 1; doodle_sprite[1][7][51] = 1; doodle_sprite[1][7][52] = 1; doodle_sprite[1][7][53] = 1; doodle_sprite[1][7][54] = 1; doodle_sprite[1][7][55] = 1; doodle_sprite[1][7][56] = 1; doodle_sprite[1][7][57] = 1; doodle_sprite[1][7][58] = 1; doodle_sprite[1][7][59] = 1; doodle_sprite[1][8][12] = 2; doodle_sprite[1][8][13] = 2; doodle_sprite[1][8][14] = 2; doodle_sprite[1][8][15] = 2; doodle_sprite[1][8][16] = 2; doodle_sprite[1][8][44] = 1; doodle_sprite[1][8][45] = 1; doodle_sprite[1][8][46] = 1; doodle_sprite[1][8][47] = 1; doodle_sprite[1][8][56] = 1; doodle_sprite[1][8][57] = 1; doodle_sprite[1][8][58] = 1; doodle_sprite[1][8][59] = 1; doodle_sprite[1][8][60] = 2; doodle_sprite[1][8][61] = 1; doodle_sprite[1][8][62] = 1; doodle_sprite[1][8][63] = 1; doodle_sprite[1][8][64] = 1; doodle_sprite[1][8][65] = 2; doodle_sprite[1][8][66] = 2; doodle_sprite[1][8][67] = 2; doodle_sprite[1][8][68] = 2; doodle_sprite[1][8][69] = 2; doodle_sprite[1][8][70] = 2; doodle_sprite[1][8][71] = 2; doodle_sprite[1][9][12] = 2; doodle_sprite[1][9][13] = 2; doodle_sprite[1][9][14] = 2; doodle_sprite[1][9][15] = 2; doodle_sprite[1][9][44] = 1; doodle_sprite[1][9][45] = 1; doodle_sprite[1][9][46] = 1; doodle_sprite[1][9][47] = 1; doodle_sprite[1][9][56] = 1; doodle_sprite[1][9][57] = 1; doodle_sprite[1][9][58] = 1; doodle_sprite[1][9][59] = 1; doodle_sprite[1][9][60] = 2; doodle_sprite[1][9][61] = 1; doodle_sprite[1][9][62] = 1; doodle_sprite[1][9][63] = 1; doodle_sprite[1][9][64] = 1; doodle_sprite[1][9][65] = 2; doodle_sprite[1][9][66] = 2; doodle_sprite[1][9][67] = 2; doodle_sprite[1][9][68] = 2; doodle_sprite[1][9][69] = 2; doodle_sprite[1][9][70] = 2; doodle_sprite[1][9][71] = 2; doodle_sprite[1][10][12] = 2; doodle_sprite[1][10][13] = 2; doodle_sprite[1][10][14] = 2; doodle_sprite[1][10][15] = 2; doodle_sprite[1][10][44] = 1; doodle_sprite[1][10][45] = 1; doodle_sprite[1][10][46] = 1; doodle_sprite[1][10][47] = 1; doodle_sprite[1][10][56] = 1; doodle_sprite[1][10][57] = 1; doodle_sprite[1][10][58] = 1; doodle_sprite[1][10][59] = 1; doodle_sprite[1][10][60] = 2; doodle_sprite[1][10][61] = 1; doodle_sprite[1][10][62] = 1; doodle_sprite[1][10][63] = 1; doodle_sprite[1][10][64] = 1; doodle_sprite[1][10][65] = 2; doodle_sprite[1][10][66] = 2; doodle_sprite[1][10][67] = 2; doodle_sprite[1][10][68] = 2; doodle_sprite[1][10][69] = 2; doodle_sprite[1][10][70] = 2; doodle_sprite[1][10][71] = 2; doodle_sprite[1][11][12] = 2; doodle_sprite[1][11][13] = 2; doodle_sprite[1][11][14] = 2; doodle_sprite[1][11][15] = 1; doodle_sprite[1][11][44] = 1; doodle_sprite[1][11][45] = 1; doodle_sprite[1][11][46] = 1; doodle_sprite[1][11][47] = 1; doodle_sprite[1][11][56] = 1; doodle_sprite[1][11][57] = 1; doodle_sprite[1][11][58] = 1; doodle_sprite[1][11][59] = 1; doodle_sprite[1][11][60] = 2; doodle_sprite[1][11][61] = 1; doodle_sprite[1][11][62] = 1; doodle_sprite[1][11][63] = 1; doodle_sprite[1][11][64] = 1; doodle_sprite[1][11][65] = 2; doodle_sprite[1][11][66] = 2; doodle_sprite[1][11][67] = 2; doodle_sprite[1][11][68] = 2; doodle_sprite[1][11][69] = 2; doodle_sprite[1][11][70] = 2; doodle_sprite[1][11][71] = 2; doodle_sprite[1][12][8] = 1; doodle_sprite[1][12][9] = 1; doodle_sprite[1][12][10] = 1; doodle_sprite[1][12][11] = 1; doodle_sprite[1][12][44] = 1; doodle_sprite[1][12][45] = 1; doodle_sprite[1][12][46] = 1; doodle_sprite[1][12][47] = 1; doodle_sprite[1][12][56] = 1; doodle_sprite[1][12][57] = 1; doodle_sprite[1][12][58] = 1; doodle_sprite[1][12][59] = 1; doodle_sprite[1][12][68] = 2; doodle_sprite[1][12][69] = 2; doodle_sprite[1][12][70] = 2; doodle_sprite[1][12][71] = 2; doodle_sprite[1][13][8] = 1; doodle_sprite[1][13][9] = 1; doodle_sprite[1][13][10] = 1; doodle_sprite[1][13][11] = 1; doodle_sprite[1][13][44] = 1; doodle_sprite[1][13][45] = 1; doodle_sprite[1][13][46] = 1; doodle_sprite[1][13][47] = 1; doodle_sprite[1][13][56] = 1; doodle_sprite[1][13][57] = 1; doodle_sprite[1][13][58] = 1; doodle_sprite[1][13][59] = 1; doodle_sprite[1][13][68] = 2; doodle_sprite[1][13][69] = 2; doodle_sprite[1][13][70] = 2; doodle_sprite[1][13][71] = 2; doodle_sprite[1][14][8] = 1; doodle_sprite[1][14][9] = 1; doodle_sprite[1][14][10] = 1; doodle_sprite[1][14][11] = 1; doodle_sprite[1][14][44] = 1; doodle_sprite[1][14][45] = 1; doodle_sprite[1][14][46] = 1; doodle_sprite[1][14][47] = 1; doodle_sprite[1][14][56] = 1; doodle_sprite[1][14][57] = 1; doodle_sprite[1][14][58] = 1; doodle_sprite[1][14][59] = 1; doodle_sprite[1][14][68] = 2; doodle_sprite[1][14][69] = 2; doodle_sprite[1][14][70] = 2; doodle_sprite[1][14][71] = 2; doodle_sprite[1][15][8] = 1; doodle_sprite[1][15][9] = 1; doodle_sprite[1][15][10] = 1; doodle_sprite[1][15][11] = 1; doodle_sprite[1][15][44] = 1; doodle_sprite[1][15][45] = 1; doodle_sprite[1][15][46] = 1; doodle_sprite[1][15][47] = 1; doodle_sprite[1][15][56] = 1; doodle_sprite[1][15][57] = 1; doodle_sprite[1][15][58] = 1; doodle_sprite[1][15][59] = 1; doodle_sprite[1][15][68] = 2; doodle_sprite[1][15][69] = 2; doodle_sprite[1][15][70] = 2; doodle_sprite[1][15][71] = 2; doodle_sprite[1][16][8] = 2; doodle_sprite[1][16][9] = 2; doodle_sprite[1][16][10] = 2; doodle_sprite[1][16][11] = 1; doodle_sprite[1][16][44] = 1; doodle_sprite[1][16][45] = 1; doodle_sprite[1][16][46] = 1; doodle_sprite[1][16][47] = 1; doodle_sprite[1][16][56] = 1; doodle_sprite[1][16][57] = 1; doodle_sprite[1][16][58] = 1; doodle_sprite[1][16][59] = 1; doodle_sprite[1][17][8] = 2; doodle_sprite[1][17][9] = 2; doodle_sprite[1][17][10] = 2; doodle_sprite[1][17][11] = 1; doodle_sprite[1][17][44] = 1; doodle_sprite[1][17][45] = 1; doodle_sprite[1][17][46] = 1; doodle_sprite[1][17][47] = 1; doodle_sprite[1][17][56] = 1; doodle_sprite[1][17][57] = 1; doodle_sprite[1][17][58] = 1; doodle_sprite[1][17][59] = 1; doodle_sprite[1][18][8] = 2; doodle_sprite[1][18][9] = 2; doodle_sprite[1][18][10] = 2; doodle_sprite[1][18][11] = 1; doodle_sprite[1][18][44] = 1; doodle_sprite[1][18][45] = 1; doodle_sprite[1][18][46] = 1; doodle_sprite[1][18][47] = 1; doodle_sprite[1][18][56] = 1; doodle_sprite[1][18][57] = 1; doodle_sprite[1][18][58] = 1; doodle_sprite[1][18][59] = 1; doodle_sprite[1][19][8] = 2; doodle_sprite[1][19][9] = 2; doodle_sprite[1][19][10] = 2; doodle_sprite[1][19][11] = 1; doodle_sprite[1][19][44] = 1; doodle_sprite[1][19][45] = 1; doodle_sprite[1][19][46] = 1; doodle_sprite[1][19][47] = 1; doodle_sprite[1][19][56] = 1; doodle_sprite[1][19][57] = 1; doodle_sprite[1][19][58] = 1; doodle_sprite[1][19][59] = 1; doodle_sprite[1][20][8] = 2; doodle_sprite[1][20][9] = 2; doodle_sprite[1][20][10] = 2; doodle_sprite[1][20][11] = 1; doodle_sprite[1][20][44] = 1; doodle_sprite[1][20][45] = 1; doodle_sprite[1][20][46] = 1; doodle_sprite[1][20][47] = 1; doodle_sprite[1][20][56] = 1; doodle_sprite[1][20][57] = 1; doodle_sprite[1][20][58] = 1; doodle_sprite[1][20][59] = 1; doodle_sprite[1][20][60] = 2; doodle_sprite[1][20][61] = 2; doodle_sprite[1][20][62] = 2; doodle_sprite[1][20][63] = 1; doodle_sprite[1][20][64] = 2; doodle_sprite[1][20][65] = 2; doodle_sprite[1][20][66] = 1; doodle_sprite[1][20][67] = 2; doodle_sprite[1][20][68] = 1; doodle_sprite[1][20][69] = 1; doodle_sprite[1][20][70] = 2; doodle_sprite[1][20][71] = 2; doodle_sprite[1][21][8] = 1; doodle_sprite[1][21][9] = 1; doodle_sprite[1][21][10] = 1; doodle_sprite[1][21][11] = 1; doodle_sprite[1][21][44] = 1; doodle_sprite[1][21][45] = 1; doodle_sprite[1][21][46] = 1; doodle_sprite[1][21][47] = 1; doodle_sprite[1][21][56] = 1; doodle_sprite[1][21][57] = 1; doodle_sprite[1][21][58] = 1; doodle_sprite[1][21][59] = 1; doodle_sprite[1][21][60] = 2; doodle_sprite[1][21][61] = 2; doodle_sprite[1][21][62] = 2; doodle_sprite[1][21][63] = 1; doodle_sprite[1][21][64] = 2; doodle_sprite[1][21][65] = 2; doodle_sprite[1][21][66] = 1; doodle_sprite[1][21][67] = 2; doodle_sprite[1][21][68] = 1; doodle_sprite[1][21][69] = 1; doodle_sprite[1][21][70] = 2; doodle_sprite[1][21][71] = 2; doodle_sprite[1][22][8] = 1; doodle_sprite[1][22][9] = 1; doodle_sprite[1][22][10] = 1; doodle_sprite[1][22][11] = 1; doodle_sprite[1][22][44] = 1; doodle_sprite[1][22][45] = 1; doodle_sprite[1][22][46] = 1; doodle_sprite[1][22][47] = 1; doodle_sprite[1][22][56] = 1; doodle_sprite[1][22][57] = 1; doodle_sprite[1][22][58] = 1; doodle_sprite[1][22][59] = 1; doodle_sprite[1][22][60] = 2; doodle_sprite[1][22][61] = 2; doodle_sprite[1][22][62] = 2; doodle_sprite[1][22][63] = 1; doodle_sprite[1][22][64] = 2; doodle_sprite[1][22][65] = 2; doodle_sprite[1][22][66] = 1; doodle_sprite[1][22][67] = 2; doodle_sprite[1][22][68] = 1; doodle_sprite[1][22][69] = 1; doodle_sprite[1][22][70] = 2; doodle_sprite[1][22][71] = 2; doodle_sprite[1][23][8] = 2; doodle_sprite[1][23][9] = 2; doodle_sprite[1][23][10] = 2; doodle_sprite[1][23][11] = 1; doodle_sprite[1][23][44] = 1; doodle_sprite[1][23][45] = 1; doodle_sprite[1][23][46] = 1; doodle_sprite[1][23][47] = 1; doodle_sprite[1][23][56] = 1; doodle_sprite[1][23][57] = 1; doodle_sprite[1][23][58] = 1; doodle_sprite[1][23][59] = 1; doodle_sprite[1][23][60] = 2; doodle_sprite[1][23][61] = 2; doodle_sprite[1][23][62] = 2; doodle_sprite[1][23][63] = 1; doodle_sprite[1][23][64] = 2; doodle_sprite[1][23][65] = 2; doodle_sprite[1][23][66] = 1; doodle_sprite[1][23][67] = 2; doodle_sprite[1][23][68] = 1; doodle_sprite[1][23][69] = 1; doodle_sprite[1][23][70] = 2; doodle_sprite[1][23][71] = 2; doodle_sprite[1][24][8] = 1; doodle_sprite[1][24][9] = 1; doodle_sprite[1][24][10] = 1; doodle_sprite[1][24][11] = 1; doodle_sprite[1][24][44] = 1; doodle_sprite[1][24][45] = 1; doodle_sprite[1][24][46] = 1; doodle_sprite[1][24][47] = 1; doodle_sprite[1][24][56] = 1; doodle_sprite[1][24][57] = 1; doodle_sprite[1][24][58] = 1; doodle_sprite[1][24][59] = 1; doodle_sprite[1][24][68] = 2; doodle_sprite[1][24][69] = 2; doodle_sprite[1][24][70] = 2; doodle_sprite[1][24][71] = 2; doodle_sprite[1][25][8] = 1; doodle_sprite[1][25][9] = 1; doodle_sprite[1][25][10] = 1; doodle_sprite[1][25][11] = 1; doodle_sprite[1][25][44] = 1; doodle_sprite[1][25][45] = 1; doodle_sprite[1][25][46] = 1; doodle_sprite[1][25][47] = 1; doodle_sprite[1][25][56] = 1; doodle_sprite[1][25][57] = 1; doodle_sprite[1][25][58] = 1; doodle_sprite[1][25][59] = 1; doodle_sprite[1][25][68] = 2; doodle_sprite[1][25][69] = 2; doodle_sprite[1][25][70] = 2; doodle_sprite[1][25][71] = 2; doodle_sprite[1][26][8] = 1; doodle_sprite[1][26][9] = 1; doodle_sprite[1][26][10] = 1; doodle_sprite[1][26][11] = 1; doodle_sprite[1][26][44] = 1; doodle_sprite[1][26][45] = 1; doodle_sprite[1][26][46] = 1; doodle_sprite[1][26][47] = 1; doodle_sprite[1][26][56] = 1; doodle_sprite[1][26][57] = 1; doodle_sprite[1][26][58] = 1; doodle_sprite[1][26][59] = 1; doodle_sprite[1][26][68] = 2; doodle_sprite[1][26][69] = 2; doodle_sprite[1][26][70] = 2; doodle_sprite[1][26][71] = 2; doodle_sprite[1][27][8] = 1; doodle_sprite[1][27][9] = 1; doodle_sprite[1][27][10] = 1; doodle_sprite[1][27][11] = 1; doodle_sprite[1][27][44] = 1; doodle_sprite[1][27][45] = 1; doodle_sprite[1][27][46] = 1; doodle_sprite[1][27][47] = 1; doodle_sprite[1][27][56] = 1; doodle_sprite[1][27][57] = 1; doodle_sprite[1][27][58] = 1; doodle_sprite[1][27][59] = 1; doodle_sprite[1][27][68] = 2; doodle_sprite[1][27][69] = 2; doodle_sprite[1][27][70] = 2; doodle_sprite[1][27][71] = 2; doodle_sprite[1][28][8] = 1; doodle_sprite[1][28][9] = 1; doodle_sprite[1][28][10] = 1; doodle_sprite[1][28][11] = 1; doodle_sprite[1][28][44] = 1; doodle_sprite[1][28][45] = 1; doodle_sprite[1][28][46] = 1; doodle_sprite[1][28][47] = 1; doodle_sprite[1][28][56] = 1; doodle_sprite[1][28][57] = 1; doodle_sprite[1][28][58] = 1; doodle_sprite[1][28][59] = 1; doodle_sprite[1][29][8] = 1; doodle_sprite[1][29][9] = 1; doodle_sprite[1][29][10] = 1; doodle_sprite[1][29][11] = 1; doodle_sprite[1][29][44] = 1; doodle_sprite[1][29][45] = 1; doodle_sprite[1][29][46] = 1; doodle_sprite[1][29][47] = 1; doodle_sprite[1][29][56] = 1; doodle_sprite[1][29][57] = 1; doodle_sprite[1][29][58] = 1; doodle_sprite[1][29][59] = 1; doodle_sprite[1][30][8] = 1; doodle_sprite[1][30][9] = 1; doodle_sprite[1][30][10] = 1; doodle_sprite[1][30][11] = 1; doodle_sprite[1][30][44] = 1; doodle_sprite[1][30][45] = 1; doodle_sprite[1][30][46] = 1; doodle_sprite[1][30][47] = 1; doodle_sprite[1][30][56] = 1; doodle_sprite[1][30][57] = 1; doodle_sprite[1][30][58] = 1; doodle_sprite[1][30][59] = 1; doodle_sprite[1][31][8] = 2; doodle_sprite[1][31][9] = 2; doodle_sprite[1][31][10] = 2; doodle_sprite[1][31][11] = 1; doodle_sprite[1][31][44] = 1; doodle_sprite[1][31][45] = 1; doodle_sprite[1][31][46] = 1; doodle_sprite[1][31][47] = 1; doodle_sprite[1][31][56] = 1; doodle_sprite[1][31][57] = 1; doodle_sprite[1][31][58] = 1; doodle_sprite[1][31][59] = 1; doodle_sprite[1][32][8] = 2; doodle_sprite[1][32][9] = 2; doodle_sprite[1][32][10] = 2; doodle_sprite[1][32][11] = 1; doodle_sprite[1][32][24] = 1; doodle_sprite[1][32][25] = 1; doodle_sprite[1][32][26] = 1; doodle_sprite[1][32][27] = 1; doodle_sprite[1][32][44] = 1; doodle_sprite[1][32][45] = 1; doodle_sprite[1][32][46] = 1; doodle_sprite[1][32][47] = 1; doodle_sprite[1][32][56] = 1; doodle_sprite[1][32][57] = 1; doodle_sprite[1][32][58] = 1; doodle_sprite[1][32][59] = 1; doodle_sprite[1][32][60] = 2; doodle_sprite[1][32][61] = 2; doodle_sprite[1][32][62] = 2; doodle_sprite[1][32][63] = 2; doodle_sprite[1][32][64] = 2; doodle_sprite[1][32][65] = 2; doodle_sprite[1][32][66] = 2; doodle_sprite[1][32][67] = 2; doodle_sprite[1][32][68] = 2; doodle_sprite[1][32][69] = 2; doodle_sprite[1][32][70] = 2; doodle_sprite[1][32][71] = 2; doodle_sprite[1][33][8] = 2; doodle_sprite[1][33][9] = 2; doodle_sprite[1][33][10] = 2; doodle_sprite[1][33][11] = 1; doodle_sprite[1][33][24] = 1; doodle_sprite[1][33][25] = 1; doodle_sprite[1][33][26] = 1; doodle_sprite[1][33][27] = 1; doodle_sprite[1][33][44] = 1; doodle_sprite[1][33][45] = 1; doodle_sprite[1][33][46] = 1; doodle_sprite[1][33][47] = 1; doodle_sprite[1][33][56] = 1; doodle_sprite[1][33][57] = 1; doodle_sprite[1][33][58] = 1; doodle_sprite[1][33][59] = 1; doodle_sprite[1][33][60] = 2; doodle_sprite[1][33][61] = 2; doodle_sprite[1][33][62] = 2; doodle_sprite[1][33][63] = 2; doodle_sprite[1][33][64] = 2; doodle_sprite[1][33][65] = 2; doodle_sprite[1][33][66] = 2; doodle_sprite[1][33][67] = 2; doodle_sprite[1][33][68] = 2; doodle_sprite[1][33][69] = 2; doodle_sprite[1][33][70] = 2; doodle_sprite[1][33][71] = 2; doodle_sprite[1][34][8] = 2; doodle_sprite[1][34][9] = 2; doodle_sprite[1][34][10] = 2; doodle_sprite[1][34][11] = 1; doodle_sprite[1][34][24] = 1; doodle_sprite[1][34][25] = 1; doodle_sprite[1][34][26] = 1; doodle_sprite[1][34][27] = 1; doodle_sprite[1][34][44] = 1; doodle_sprite[1][34][45] = 1; doodle_sprite[1][34][46] = 1; doodle_sprite[1][34][47] = 1; doodle_sprite[1][34][56] = 1; doodle_sprite[1][34][57] = 1; doodle_sprite[1][34][58] = 1; doodle_sprite[1][34][59] = 1; doodle_sprite[1][34][60] = 2; doodle_sprite[1][34][61] = 2; doodle_sprite[1][34][62] = 2; doodle_sprite[1][34][63] = 2; doodle_sprite[1][34][64] = 2; doodle_sprite[1][34][65] = 2; doodle_sprite[1][34][66] = 2; doodle_sprite[1][34][67] = 2; doodle_sprite[1][34][68] = 2; doodle_sprite[1][34][69] = 2; doodle_sprite[1][34][70] = 2; doodle_sprite[1][34][71] = 2; doodle_sprite[1][35][8] = 2; doodle_sprite[1][35][9] = 2; doodle_sprite[1][35][10] = 2; doodle_sprite[1][35][11] = 1; doodle_sprite[1][35][24] = 1; doodle_sprite[1][35][25] = 1; doodle_sprite[1][35][26] = 1; doodle_sprite[1][35][27] = 1; doodle_sprite[1][35][44] = 1; doodle_sprite[1][35][45] = 1; doodle_sprite[1][35][46] = 1; doodle_sprite[1][35][47] = 1; doodle_sprite[1][35][56] = 1; doodle_sprite[1][35][57] = 1; doodle_sprite[1][35][58] = 1; doodle_sprite[1][35][59] = 1; doodle_sprite[1][35][60] = 2; doodle_sprite[1][35][61] = 2; doodle_sprite[1][35][62] = 2; doodle_sprite[1][35][63] = 2; doodle_sprite[1][35][64] = 2; doodle_sprite[1][35][65] = 2; doodle_sprite[1][35][66] = 2; doodle_sprite[1][35][67] = 2; doodle_sprite[1][35][68] = 2; doodle_sprite[1][35][69] = 2; doodle_sprite[1][35][70] = 2; doodle_sprite[1][35][71] = 2; doodle_sprite[1][36][8] = 2; doodle_sprite[1][36][9] = 2; doodle_sprite[1][36][10] = 2; doodle_sprite[1][36][11] = 1; doodle_sprite[1][36][44] = 1; doodle_sprite[1][36][45] = 1; doodle_sprite[1][36][46] = 1; doodle_sprite[1][36][47] = 1; doodle_sprite[1][36][56] = 1; doodle_sprite[1][36][57] = 1; doodle_sprite[1][36][58] = 1; doodle_sprite[1][36][59] = 1; doodle_sprite[1][36][68] = 2; doodle_sprite[1][36][69] = 2; doodle_sprite[1][36][70] = 2; doodle_sprite[1][36][71] = 2; doodle_sprite[1][37][8] = 2; doodle_sprite[1][37][9] = 2; doodle_sprite[1][37][10] = 2; doodle_sprite[1][37][11] = 1; doodle_sprite[1][37][44] = 1; doodle_sprite[1][37][45] = 1; doodle_sprite[1][37][46] = 1; doodle_sprite[1][37][47] = 1; doodle_sprite[1][37][56] = 1; doodle_sprite[1][37][57] = 1; doodle_sprite[1][37][58] = 1; doodle_sprite[1][37][59] = 1; doodle_sprite[1][37][68] = 2; doodle_sprite[1][37][69] = 2; doodle_sprite[1][37][70] = 2; doodle_sprite[1][37][71] = 2; doodle_sprite[1][38][8] = 2; doodle_sprite[1][38][9] = 2; doodle_sprite[1][38][10] = 2; doodle_sprite[1][38][11] = 2; doodle_sprite[1][38][44] = 1; doodle_sprite[1][38][45] = 1; doodle_sprite[1][38][46] = 1; doodle_sprite[1][38][47] = 1; doodle_sprite[1][38][56] = 1; doodle_sprite[1][38][57] = 1; doodle_sprite[1][38][58] = 1; doodle_sprite[1][38][59] = 1; doodle_sprite[1][38][68] = 2; doodle_sprite[1][38][69] = 2; doodle_sprite[1][38][70] = 2; doodle_sprite[1][38][71] = 2; doodle_sprite[1][39][8] = 2; doodle_sprite[1][39][9] = 2; doodle_sprite[1][39][10] = 2; doodle_sprite[1][39][11] = 2; doodle_sprite[1][39][44] = 1; doodle_sprite[1][39][45] = 1; doodle_sprite[1][39][46] = 1; doodle_sprite[1][39][47] = 1; doodle_sprite[1][39][56] = 1; doodle_sprite[1][39][57] = 1; doodle_sprite[1][39][58] = 1; doodle_sprite[1][39][59] = 1; doodle_sprite[1][39][68] = 2; doodle_sprite[1][39][69] = 2; doodle_sprite[1][39][70] = 2; doodle_sprite[1][39][71] = 2; doodle_sprite[1][40][8] = 2; doodle_sprite[1][40][9] = 2; doodle_sprite[1][40][10] = 2; doodle_sprite[1][40][11] = 2; doodle_sprite[1][40][24] = 1; doodle_sprite[1][40][25] = 1; doodle_sprite[1][40][26] = 1; doodle_sprite[1][40][27] = 1; doodle_sprite[1][40][44] = 1; doodle_sprite[1][40][45] = 1; doodle_sprite[1][40][46] = 1; doodle_sprite[1][40][47] = 1; doodle_sprite[1][40][56] = 1; doodle_sprite[1][40][57] = 1; doodle_sprite[1][40][58] = 1; doodle_sprite[1][40][59] = 1; doodle_sprite[1][41][8] = 2; doodle_sprite[1][41][9] = 2; doodle_sprite[1][41][10] = 2; doodle_sprite[1][41][11] = 2; doodle_sprite[1][41][24] = 1; doodle_sprite[1][41][25] = 1; doodle_sprite[1][41][26] = 1; doodle_sprite[1][41][27] = 1; doodle_sprite[1][41][44] = 1; doodle_sprite[1][41][45] = 1; doodle_sprite[1][41][46] = 1; doodle_sprite[1][41][47] = 1; doodle_sprite[1][41][56] = 1; doodle_sprite[1][41][57] = 1; doodle_sprite[1][41][58] = 1; doodle_sprite[1][41][59] = 1; doodle_sprite[1][42][8] = 2; doodle_sprite[1][42][9] = 2; doodle_sprite[1][42][10] = 2; doodle_sprite[1][42][11] = 2; doodle_sprite[1][42][24] = 1; doodle_sprite[1][42][25] = 1; doodle_sprite[1][42][26] = 1; doodle_sprite[1][42][27] = 1; doodle_sprite[1][42][44] = 1; doodle_sprite[1][42][45] = 1; doodle_sprite[1][42][46] = 1; doodle_sprite[1][42][47] = 1; doodle_sprite[1][42][56] = 1; doodle_sprite[1][42][57] = 1; doodle_sprite[1][42][58] = 1; doodle_sprite[1][42][59] = 1; doodle_sprite[1][43][8] = 2; doodle_sprite[1][43][9] = 2; doodle_sprite[1][43][10] = 2; doodle_sprite[1][43][11] = 2; doodle_sprite[1][43][24] = 1; doodle_sprite[1][43][25] = 1; doodle_sprite[1][43][26] = 1; doodle_sprite[1][43][27] = 1; doodle_sprite[1][43][44] = 1; doodle_sprite[1][43][45] = 1; doodle_sprite[1][43][46] = 1; doodle_sprite[1][43][47] = 1; doodle_sprite[1][43][56] = 1; doodle_sprite[1][43][57] = 1; doodle_sprite[1][43][58] = 1; doodle_sprite[1][43][59] = 1; doodle_sprite[1][44][12] = 2; doodle_sprite[1][44][13] = 2; doodle_sprite[1][44][14] = 2; doodle_sprite[1][44][15] = 2; doodle_sprite[1][44][16] = 2; doodle_sprite[1][44][44] = 1; doodle_sprite[1][44][45] = 1; doodle_sprite[1][44][46] = 1; doodle_sprite[1][44][47] = 1; doodle_sprite[1][44][56] = 1; doodle_sprite[1][44][57] = 1; doodle_sprite[1][44][58] = 1; doodle_sprite[1][44][59] = 1; doodle_sprite[1][44][60] = 2; doodle_sprite[1][44][61] = 2; doodle_sprite[1][44][62] = 2; doodle_sprite[1][44][63] = 2; doodle_sprite[1][44][64] = 2; doodle_sprite[1][44][65] = 2; doodle_sprite[1][44][66] = 2; doodle_sprite[1][44][67] = 2; doodle_sprite[1][44][68] = 2; doodle_sprite[1][44][69] = 2; doodle_sprite[1][44][70] = 2; doodle_sprite[1][44][71] = 2; doodle_sprite[1][45][12] = 2; doodle_sprite[1][45][13] = 2; doodle_sprite[1][45][14] = 2; doodle_sprite[1][45][15] = 2; doodle_sprite[1][45][16] = 2; doodle_sprite[1][45][44] = 1; doodle_sprite[1][45][45] = 1; doodle_sprite[1][45][46] = 1; doodle_sprite[1][45][47] = 1; doodle_sprite[1][45][56] = 1; doodle_sprite[1][45][57] = 1; doodle_sprite[1][45][58] = 1; doodle_sprite[1][45][59] = 1; doodle_sprite[1][45][60] = 2; doodle_sprite[1][45][61] = 2; doodle_sprite[1][45][62] = 2; doodle_sprite[1][45][63] = 2; doodle_sprite[1][45][64] = 2; doodle_sprite[1][45][65] = 2; doodle_sprite[1][45][66] = 2; doodle_sprite[1][45][67] = 2; doodle_sprite[1][45][68] = 2; doodle_sprite[1][45][69] = 2; doodle_sprite[1][45][70] = 2; doodle_sprite[1][45][71] = 2; doodle_sprite[1][46][12] = 2; doodle_sprite[1][46][13] = 2; doodle_sprite[1][46][14] = 2; doodle_sprite[1][46][15] = 2; doodle_sprite[1][46][16] = 2; doodle_sprite[1][46][44] = 1; doodle_sprite[1][46][45] = 1; doodle_sprite[1][46][46] = 1; doodle_sprite[1][46][47] = 1; doodle_sprite[1][46][56] = 1; doodle_sprite[1][46][57] = 1; doodle_sprite[1][46][58] = 1; doodle_sprite[1][46][59] = 1; doodle_sprite[1][46][60] = 2; doodle_sprite[1][46][61] = 2; doodle_sprite[1][46][62] = 2; doodle_sprite[1][46][63] = 2; doodle_sprite[1][46][64] = 2; doodle_sprite[1][46][65] = 2; doodle_sprite[1][46][66] = 2; doodle_sprite[1][46][67] = 2; doodle_sprite[1][46][68] = 2; doodle_sprite[1][46][69] = 2; doodle_sprite[1][46][70] = 2; doodle_sprite[1][46][71] = 2; doodle_sprite[1][47][12] = 2; doodle_sprite[1][47][13] = 2; doodle_sprite[1][47][14] = 2; doodle_sprite[1][47][15] = 2; doodle_sprite[1][47][16] = 2; doodle_sprite[1][47][44] = 1; doodle_sprite[1][47][45] = 1; doodle_sprite[1][47][46] = 1; doodle_sprite[1][47][47] = 1; doodle_sprite[1][47][56] = 1; doodle_sprite[1][47][57] = 1; doodle_sprite[1][47][58] = 1; doodle_sprite[1][47][59] = 1; doodle_sprite[1][47][60] = 2; doodle_sprite[1][47][61] = 2; doodle_sprite[1][47][62] = 2; doodle_sprite[1][47][63] = 2; doodle_sprite[1][47][64] = 2; doodle_sprite[1][47][65] = 2; doodle_sprite[1][47][66] = 2; doodle_sprite[1][47][67] = 2; doodle_sprite[1][47][68] = 2; doodle_sprite[1][47][69] = 2; doodle_sprite[1][47][70] = 2; doodle_sprite[1][47][71] = 2; doodle_sprite[1][48][16] = 2; doodle_sprite[1][48][17] = 2; doodle_sprite[1][48][18] = 2; doodle_sprite[1][48][19] = 2; doodle_sprite[1][48][20] = 2; doodle_sprite[1][48][21] = 2; doodle_sprite[1][48][22] = 2; doodle_sprite[1][48][23] = 2; doodle_sprite[1][48][24] = 2; doodle_sprite[1][48][25] = 2; doodle_sprite[1][48][26] = 2; doodle_sprite[1][48][27] = 1; doodle_sprite[1][48][36] = 1; doodle_sprite[1][48][37] = 1; doodle_sprite[1][48][38] = 1; doodle_sprite[1][48][39] = 1; doodle_sprite[1][48][40] = 1; doodle_sprite[1][48][41] = 1; doodle_sprite[1][48][42] = 1; doodle_sprite[1][48][43] = 1; doodle_sprite[1][48][44] = 1; doodle_sprite[1][48][45] = 1; doodle_sprite[1][48][46] = 1; doodle_sprite[1][48][47] = 1; doodle_sprite[1][48][48] = 1; doodle_sprite[1][48][49] = 1; doodle_sprite[1][48][50] = 1; doodle_sprite[1][48][51] = 1; doodle_sprite[1][48][52] = 1; doodle_sprite[1][48][53] = 1; doodle_sprite[1][48][54] = 1; doodle_sprite[1][48][55] = 1; doodle_sprite[1][48][56] = 1; doodle_sprite[1][48][57] = 1; doodle_sprite[1][48][58] = 1; doodle_sprite[1][48][59] = 1; doodle_sprite[1][48][68] = 2; doodle_sprite[1][48][69] = 2; doodle_sprite[1][48][70] = 2; doodle_sprite[1][48][71] = 2; doodle_sprite[1][49][16] = 2; doodle_sprite[1][49][17] = 2; doodle_sprite[1][49][18] = 2; doodle_sprite[1][49][19] = 2; doodle_sprite[1][49][20] = 2; doodle_sprite[1][49][21] = 2; doodle_sprite[1][49][22] = 2; doodle_sprite[1][49][23] = 2; doodle_sprite[1][49][24] = 1; doodle_sprite[1][49][25] = 1; doodle_sprite[1][49][26] = 1; doodle_sprite[1][49][27] = 1; doodle_sprite[1][49][36] = 1; doodle_sprite[1][49][37] = 1; doodle_sprite[1][49][38] = 1; doodle_sprite[1][49][39] = 1; doodle_sprite[1][49][40] = 1; doodle_sprite[1][49][41] = 1; doodle_sprite[1][49][42] = 1; doodle_sprite[1][49][43] = 1; doodle_sprite[1][49][44] = 1; doodle_sprite[1][49][45] = 1; doodle_sprite[1][49][46] = 1; doodle_sprite[1][49][47] = 1; doodle_sprite[1][49][48] = 1; doodle_sprite[1][49][49] = 1; doodle_sprite[1][49][50] = 1; doodle_sprite[1][49][51] = 1; doodle_sprite[1][49][52] = 1; doodle_sprite[1][49][53] = 1; doodle_sprite[1][49][54] = 1; doodle_sprite[1][49][55] = 1; doodle_sprite[1][49][56] = 1; doodle_sprite[1][49][57] = 1; doodle_sprite[1][49][58] = 1; doodle_sprite[1][49][59] = 1; doodle_sprite[1][49][68] = 2; doodle_sprite[1][49][69] = 2; doodle_sprite[1][49][70] = 2; doodle_sprite[1][49][71] = 2; doodle_sprite[1][50][16] = 2; doodle_sprite[1][50][17] = 2; doodle_sprite[1][50][18] = 2; doodle_sprite[1][50][19] = 2; doodle_sprite[1][50][20] = 2; doodle_sprite[1][50][21] = 2; doodle_sprite[1][50][22] = 2; doodle_sprite[1][50][23] = 2; doodle_sprite[1][50][24] = 1; doodle_sprite[1][50][25] = 1; doodle_sprite[1][50][26] = 1; doodle_sprite[1][50][27] = 1; doodle_sprite[1][50][36] = 1; doodle_sprite[1][50][37] = 1; doodle_sprite[1][50][38] = 1; doodle_sprite[1][50][39] = 1; doodle_sprite[1][50][40] = 1; doodle_sprite[1][50][41] = 1; doodle_sprite[1][50][42] = 1; doodle_sprite[1][50][43] = 1; doodle_sprite[1][50][44] = 1; doodle_sprite[1][50][45] = 1; doodle_sprite[1][50][46] = 1; doodle_sprite[1][50][47] = 1; doodle_sprite[1][50][48] = 1; doodle_sprite[1][50][49] = 1; doodle_sprite[1][50][50] = 1; doodle_sprite[1][50][51] = 1; doodle_sprite[1][50][52] = 1; doodle_sprite[1][50][53] = 1; doodle_sprite[1][50][54] = 1; doodle_sprite[1][50][55] = 1; doodle_sprite[1][50][56] = 1; doodle_sprite[1][50][57] = 2; doodle_sprite[1][50][58] = 2; doodle_sprite[1][50][59] = 2; doodle_sprite[1][50][68] = 2; doodle_sprite[1][50][69] = 2; doodle_sprite[1][50][70] = 2; doodle_sprite[1][50][71] = 2; doodle_sprite[1][51][16] = 2; doodle_sprite[1][51][17] = 2; doodle_sprite[1][51][18] = 2; doodle_sprite[1][51][19] = 2; doodle_sprite[1][51][20] = 2; doodle_sprite[1][51][21] = 2; doodle_sprite[1][51][22] = 2; doodle_sprite[1][51][23] = 2; doodle_sprite[1][51][24] = 1; doodle_sprite[1][51][25] = 1; doodle_sprite[1][51][26] = 1; doodle_sprite[1][51][27] = 1; doodle_sprite[1][51][35] = 2; doodle_sprite[1][51][36] = 1; doodle_sprite[1][51][37] = 1; doodle_sprite[1][51][38] = 1; doodle_sprite[1][51][39] = 1; doodle_sprite[1][51][40] = 1; doodle_sprite[1][51][41] = 1; doodle_sprite[1][51][42] = 1; doodle_sprite[1][51][43] = 1; doodle_sprite[1][51][44] = 1; doodle_sprite[1][51][45] = 1; doodle_sprite[1][51][46] = 1; doodle_sprite[1][51][47] = 1; doodle_sprite[1][51][48] = 1; doodle_sprite[1][51][49] = 1; doodle_sprite[1][51][50] = 1; doodle_sprite[1][51][51] = 1; doodle_sprite[1][51][52] = 1; doodle_sprite[1][51][53] = 1; doodle_sprite[1][51][54] = 1; doodle_sprite[1][51][55] = 1; doodle_sprite[1][51][56] = 1; doodle_sprite[1][51][57] = 2; doodle_sprite[1][51][58] = 2; doodle_sprite[1][51][59] = 2; doodle_sprite[1][51][68] = 2; doodle_sprite[1][51][69] = 2; doodle_sprite[1][51][70] = 2; doodle_sprite[1][51][71] = 2; doodle_sprite[1][52][24] = 1; doodle_sprite[1][52][25] = 1; doodle_sprite[1][52][26] = 1; doodle_sprite[1][52][27] = 1; doodle_sprite[1][52][32] = 1; doodle_sprite[1][52][33] = 1; doodle_sprite[1][52][34] = 1; doodle_sprite[1][52][35] = 1; doodle_sprite[1][53][24] = 1; doodle_sprite[1][53][25] = 1; doodle_sprite[1][53][26] = 1; doodle_sprite[1][53][27] = 1; doodle_sprite[1][53][32] = 1; doodle_sprite[1][53][33] = 1; doodle_sprite[1][53][34] = 1; doodle_sprite[1][53][35] = 1; doodle_sprite[1][54][24] = 1; doodle_sprite[1][54][25] = 1; doodle_sprite[1][54][26] = 1; doodle_sprite[1][54][27] = 1; doodle_sprite[1][54][32] = 1; doodle_sprite[1][54][33] = 1; doodle_sprite[1][54][34] = 1; doodle_sprite[1][54][35] = 1; doodle_sprite[1][55][24] = 1; doodle_sprite[1][55][25] = 1; doodle_sprite[1][55][26] = 1; doodle_sprite[1][55][27] = 1; doodle_sprite[1][55][32] = 1; doodle_sprite[1][55][33] = 1; doodle_sprite[1][55][34] = 1; doodle_sprite[1][55][35] = 1; doodle_sprite[1][56][24] = 1; doodle_sprite[1][56][25] = 1; doodle_sprite[1][56][26] = 1; doodle_sprite[1][56][27] = 1; doodle_sprite[1][56][32] = 1; doodle_sprite[1][56][33] = 1; doodle_sprite[1][56][34] = 1; doodle_sprite[1][56][35] = 1; doodle_sprite[1][57][24] = 1; doodle_sprite[1][57][25] = 1; doodle_sprite[1][57][26] = 1; doodle_sprite[1][57][27] = 1; doodle_sprite[1][57][32] = 1; doodle_sprite[1][57][33] = 1; doodle_sprite[1][57][34] = 1; doodle_sprite[1][57][35] = 1; doodle_sprite[1][58][24] = 1; doodle_sprite[1][58][25] = 1; doodle_sprite[1][58][26] = 1; doodle_sprite[1][58][27] = 1; doodle_sprite[1][58][32] = 1; doodle_sprite[1][58][33] = 1; doodle_sprite[1][58][34] = 1; doodle_sprite[1][58][35] = 1; doodle_sprite[1][59][24] = 1; doodle_sprite[1][59][25] = 1; doodle_sprite[1][59][26] = 1; doodle_sprite[1][59][27] = 1; doodle_sprite[1][59][32] = 1; doodle_sprite[1][59][33] = 1; doodle_sprite[1][59][34] = 1; doodle_sprite[1][59][35] = 1; doodle_sprite[1][60][24] = 1; doodle_sprite[1][60][25] = 1; doodle_sprite[1][60][26] = 1; doodle_sprite[1][60][27] = 1; doodle_sprite[1][60][32] = 1; doodle_sprite[1][60][33] = 1; doodle_sprite[1][60][34] = 1; doodle_sprite[1][60][35] = 1; doodle_sprite[1][61][24] = 1; doodle_sprite[1][61][25] = 1; doodle_sprite[1][61][26] = 1; doodle_sprite[1][61][27] = 1; doodle_sprite[1][61][32] = 1; doodle_sprite[1][61][33] = 1; doodle_sprite[1][61][34] = 1; doodle_sprite[1][61][35] = 1; doodle_sprite[1][62][24] = 1; doodle_sprite[1][62][25] = 1; doodle_sprite[1][62][26] = 1; doodle_sprite[1][62][27] = 1; doodle_sprite[1][62][32] = 1; doodle_sprite[1][62][33] = 1; doodle_sprite[1][62][34] = 1; doodle_sprite[1][62][35] = 1; doodle_sprite[1][63][24] = 1; doodle_sprite[1][63][25] = 1; doodle_sprite[1][63][26] = 1; doodle_sprite[1][63][27] = 1; doodle_sprite[1][63][32] = 1; doodle_sprite[1][63][33] = 1; doodle_sprite[1][63][34] = 1; doodle_sprite[1][63][35] = 1; doodle_sprite[1][64][24] = 1; doodle_sprite[1][64][25] = 1; doodle_sprite[1][64][26] = 1; doodle_sprite[1][64][27] = 1; doodle_sprite[1][64][28] = 1; doodle_sprite[1][64][29] = 1; doodle_sprite[1][64][30] = 1; doodle_sprite[1][64][31] = 1; doodle_sprite[1][64][32] = 1; doodle_sprite[1][64][33] = 1; doodle_sprite[1][64][34] = 1; doodle_sprite[1][64][35] = 1; doodle_sprite[1][65][24] = 1; doodle_sprite[1][65][25] = 1; doodle_sprite[1][65][26] = 1; doodle_sprite[1][65][27] = 1; doodle_sprite[1][65][28] = 1; doodle_sprite[1][65][29] = 1; doodle_sprite[1][65][30] = 1; doodle_sprite[1][65][31] = 1; doodle_sprite[1][65][32] = 1; doodle_sprite[1][65][33] = 1; doodle_sprite[1][65][34] = 1; doodle_sprite[1][65][35] = 1; doodle_sprite[1][66][24] = 1; doodle_sprite[1][66][25] = 1; doodle_sprite[1][66][26] = 1; doodle_sprite[1][66][27] = 1; doodle_sprite[1][66][28] = 1; doodle_sprite[1][66][29] = 1; doodle_sprite[1][66][30] = 1; doodle_sprite[1][66][31] = 1; doodle_sprite[1][66][32] = 1; doodle_sprite[1][66][33] = 1; doodle_sprite[1][66][34] = 1; doodle_sprite[1][66][35] = 1; doodle_sprite[1][67][24] = 1; doodle_sprite[1][67][25] = 1; doodle_sprite[1][67][26] = 1; doodle_sprite[1][67][27] = 1; doodle_sprite[1][67][28] = 1; doodle_sprite[1][67][29] = 1; doodle_sprite[1][67][30] = 1; doodle_sprite[1][67][31] = 1; doodle_sprite[1][67][32] = 1; doodle_sprite[1][67][33] = 1; doodle_sprite[1][67][34] = 1; doodle_sprite[1][67][35] = 1; doodle_sprite[1][68][24] = 2; doodle_sprite[1][68][25] = 2; doodle_sprite[1][68][26] = 2; doodle_sprite[1][68][27] = 1; doodle_sprite[1][68][32] = 1; doodle_sprite[1][68][33] = 1; doodle_sprite[1][68][34] = 1; doodle_sprite[1][68][35] = 1; doodle_sprite[1][69][24] = 2; doodle_sprite[1][69][25] = 2; doodle_sprite[1][69][26] = 2; doodle_sprite[1][69][27] = 1; doodle_sprite[1][69][32] = 1; doodle_sprite[1][69][33] = 1; doodle_sprite[1][69][34] = 1; doodle_sprite[1][69][35] = 1; doodle_sprite[1][70][24] = 2; doodle_sprite[1][70][25] = 2; doodle_sprite[1][70][26] = 2; doodle_sprite[1][70][27] = 1; doodle_sprite[1][70][32] = 1; doodle_sprite[1][70][33] = 1; doodle_sprite[1][70][34] = 1; doodle_sprite[1][70][35] = 1; doodle_sprite[1][71][24] = 2; doodle_sprite[1][71][25] = 2; doodle_sprite[1][71][26] = 2; doodle_sprite[1][71][27] = 1; doodle_sprite[1][71][32] = 1; doodle_sprite[1][71][33] = 1; doodle_sprite[1][71][34] = 1; doodle_sprite[1][71][35] = 1; doodle_sprite[1][72][24] = 2; doodle_sprite[1][72][25] = 2; doodle_sprite[1][72][26] = 2; doodle_sprite[1][72][27] = 1; doodle_sprite[1][72][28] = 1; doodle_sprite[1][72][29] = 1; doodle_sprite[1][72][30] = 1; doodle_sprite[1][72][31] = 1; doodle_sprite[1][72][32] = 1; doodle_sprite[1][72][33] = 2; doodle_sprite[1][72][34] = 2; doodle_sprite[1][72][35] = 2; doodle_sprite[1][73][24] = 2; doodle_sprite[1][73][25] = 2; doodle_sprite[1][73][26] = 2; doodle_sprite[1][73][27] = 2; doodle_sprite[1][73][28] = 2; doodle_sprite[1][73][29] = 2; doodle_sprite[1][73][30] = 2; doodle_sprite[1][73][31] = 2; doodle_sprite[1][73][32] = 2; doodle_sprite[1][73][33] = 2; doodle_sprite[1][73][34] = 2; doodle_sprite[1][73][35] = 2; doodle_sprite[1][74][24] = 2; doodle_sprite[1][74][25] = 2; doodle_sprite[1][74][26] = 2; doodle_sprite[1][74][27] = 2; doodle_sprite[1][74][28] = 2; doodle_sprite[1][74][29] = 2; doodle_sprite[1][74][30] = 2; doodle_sprite[1][74][31] = 2; doodle_sprite[1][74][32] = 2; doodle_sprite[1][74][33] = 2; doodle_sprite[1][74][34] = 2; doodle_sprite[1][74][35] = 2; doodle_sprite[1][75][24] = 2; doodle_sprite[1][75][25] = 2; doodle_sprite[1][75][26] = 2; doodle_sprite[1][75][27] = 2; doodle_sprite[1][75][28] = 2; doodle_sprite[1][75][29] = 2; doodle_sprite[1][75][30] = 2; doodle_sprite[1][75][31] = 2; doodle_sprite[1][75][32] = 2; doodle_sprite[1][75][33] = 2; doodle_sprite[1][75][34] = 2; doodle_sprite[1][75][35] = 2;
					platform_sprite[0][5][10] = 1; platform_sprite[0][5][11] = 1; platform_sprite[0][5][12] = 1; platform_sprite[0][5][13] = 1; platform_sprite[0][5][14] = 1; platform_sprite[0][5][15] = 1; platform_sprite[0][5][16] = 1; platform_sprite[0][5][17] = 1; platform_sprite[0][5][18] = 1; platform_sprite[0][5][19] = 1; platform_sprite[0][6][10] = 1; platform_sprite[0][6][11] = 1; platform_sprite[0][6][12] = 1; platform_sprite[0][6][13] = 1; platform_sprite[0][6][14] = 1; platform_sprite[0][6][15] = 1; platform_sprite[0][6][16] = 1; platform_sprite[0][6][17] = 1; platform_sprite[0][6][18] = 1; platform_sprite[0][6][19] = 1; platform_sprite[0][7][10] = 1; platform_sprite[0][7][11] = 1; platform_sprite[0][7][12] = 1; platform_sprite[0][7][13] = 1; platform_sprite[0][7][14] = 1; platform_sprite[0][7][15] = 1; platform_sprite[0][7][16] = 1; platform_sprite[0][7][17] = 1; platform_sprite[0][7][18] = 1; platform_sprite[0][7][19] = 1; platform_sprite[0][8][10] = 1; platform_sprite[0][8][11] = 1; platform_sprite[0][8][12] = 1; platform_sprite[0][8][13] = 1; platform_sprite[0][8][14] = 1; platform_sprite[0][8][15] = 1; platform_sprite[0][8][16] = 1; platform_sprite[0][8][17] = 1; platform_sprite[0][8][18] = 1; platform_sprite[0][8][19] = 1; platform_sprite[0][9][10] = 1; platform_sprite[0][9][11] = 1; platform_sprite[0][9][12] = 1; platform_sprite[0][9][13] = 1; platform_sprite[0][9][14] = 1; platform_sprite[0][9][15] = 1; platform_sprite[0][9][16] = 1; platform_sprite[0][9][17] = 1; platform_sprite[0][9][18] = 1; platform_sprite[0][9][19] = 1; platform_sprite[0][9][20] = 1; platform_sprite[0][9][21] = 1; platform_sprite[0][9][22] = 1; platform_sprite[0][9][23] = 1; platform_sprite[0][9][24] = 1; platform_sprite[0][10][5] = 1; platform_sprite[0][10][6] = 1; platform_sprite[0][10][7] = 1; platform_sprite[0][10][8] = 1; platform_sprite[0][10][9] = 1; platform_sprite[0][10][20] = 1; platform_sprite[0][10][21] = 1; platform_sprite[0][10][22] = 1; platform_sprite[0][10][23] = 1; platform_sprite[0][10][24] = 1; platform_sprite[0][11][5] = 1; platform_sprite[0][11][6] = 1; platform_sprite[0][11][7] = 1; platform_sprite[0][11][8] = 1; platform_sprite[0][11][9] = 1; platform_sprite[0][11][20] = 1; platform_sprite[0][11][21] = 1; platform_sprite[0][11][22] = 1; platform_sprite[0][11][23] = 1; platform_sprite[0][11][24] = 1; platform_sprite[0][12][5] = 1; platform_sprite[0][12][6] = 1; platform_sprite[0][12][7] = 1; platform_sprite[0][12][8] = 1; platform_sprite[0][12][9] = 1; platform_sprite[0][12][20] = 1; platform_sprite[0][12][21] = 1; platform_sprite[0][12][22] = 1; platform_sprite[0][12][23] = 1; platform_sprite[0][12][24] = 1; platform_sprite[0][13][5] = 1; platform_sprite[0][13][6] = 1; platform_sprite[0][13][7] = 1; platform_sprite[0][13][8] = 1; platform_sprite[0][13][9] = 1; platform_sprite[0][13][20] = 1; platform_sprite[0][13][21] = 1; platform_sprite[0][13][22] = 1; platform_sprite[0][13][23] = 1; platform_sprite[0][13][24] = 1; platform_sprite[0][14][5] = 1; platform_sprite[0][14][6] = 1; platform_sprite[0][14][7] = 1; platform_sprite[0][14][8] = 1; platform_sprite[0][14][9] = 1; platform_sprite[0][14][20] = 1; platform_sprite[0][14][21] = 1; platform_sprite[0][14][22] = 1; platform_sprite[0][14][23] = 1; platform_sprite[0][14][24] = 1; platform_sprite[0][15][5] = 1; platform_sprite[0][15][6] = 1; platform_sprite[0][15][7] = 1; platform_sprite[0][15][8] = 1; platform_sprite[0][15][9] = 1; platform_sprite[0][15][20] = 1; platform_sprite[0][15][21] = 1; platform_sprite[0][15][22] = 1; platform_sprite[0][15][23] = 1; platform_sprite[0][15][24] = 1; platform_sprite[0][16][5] = 1; platform_sprite[0][16][6] = 1; platform_sprite[0][16][7] = 1; platform_sprite[0][16][8] = 1; platform_sprite[0][16][9] = 1; platform_sprite[0][16][20] = 1; platform_sprite[0][16][21] = 1; platform_sprite[0][16][22] = 1; platform_sprite[0][16][23] = 1; platform_sprite[0][16][24] = 1; platform_sprite[0][17][5] = 1; platform_sprite[0][17][6] = 1; platform_sprite[0][17][7] = 1; platform_sprite[0][17][8] = 1; platform_sprite[0][17][9] = 1; platform_sprite[0][17][20] = 1; platform_sprite[0][17][21] = 1; platform_sprite[0][17][22] = 1; platform_sprite[0][17][23] = 1; platform_sprite[0][17][24] = 1; platform_sprite[0][18][5] = 1; platform_sprite[0][18][6] = 1; platform_sprite[0][18][7] = 1; platform_sprite[0][18][8] = 1; platform_sprite[0][18][9] = 1; platform_sprite[0][18][20] = 1; platform_sprite[0][18][21] = 1; platform_sprite[0][18][22] = 1; platform_sprite[0][18][23] = 1; platform_sprite[0][18][24] = 1; platform_sprite[0][19][5] = 1; platform_sprite[0][19][6] = 1; platform_sprite[0][19][7] = 1; platform_sprite[0][19][8] = 1; platform_sprite[0][19][9] = 1; platform_sprite[0][19][20] = 1; platform_sprite[0][19][21] = 1; platform_sprite[0][19][22] = 1; platform_sprite[0][19][23] = 1; platform_sprite[0][19][24] = 1; platform_sprite[0][20][5] = 1; platform_sprite[0][20][6] = 1; platform_sprite[0][20][7] = 1; platform_sprite[0][20][8] = 1; platform_sprite[0][20][9] = 1; platform_sprite[0][20][20] = 1; platform_sprite[0][20][21] = 1; platform_sprite[0][20][22] = 1; platform_sprite[0][20][23] = 1; platform_sprite[0][20][24] = 1; platform_sprite[0][21][5] = 1; platform_sprite[0][21][6] = 1; platform_sprite[0][21][7] = 1; platform_sprite[0][21][8] = 1; platform_sprite[0][21][9] = 1; platform_sprite[0][21][20] = 1; platform_sprite[0][21][21] = 1; platform_sprite[0][21][22] = 1; platform_sprite[0][21][23] = 1; platform_sprite[0][21][24] = 1; platform_sprite[0][22][5] = 1; platform_sprite[0][22][6] = 1; platform_sprite[0][22][7] = 1; platform_sprite[0][22][8] = 1; platform_sprite[0][22][9] = 1; platform_sprite[0][22][20] = 1; platform_sprite[0][22][21] = 1; platform_sprite[0][22][22] = 1; platform_sprite[0][22][23] = 1; platform_sprite[0][22][24] = 1; platform_sprite[0][23][5] = 1; platform_sprite[0][23][6] = 1; platform_sprite[0][23][7] = 1; platform_sprite[0][23][8] = 1; platform_sprite[0][23][9] = 1; platform_sprite[0][23][20] = 1; platform_sprite[0][23][21] = 1; platform_sprite[0][23][22] = 1; platform_sprite[0][23][23] = 1; platform_sprite[0][23][24] = 1; platform_sprite[0][24][5] = 1; platform_sprite[0][24][6] = 1; platform_sprite[0][24][7] = 1; platform_sprite[0][24][8] = 1; platform_sprite[0][24][9] = 1; platform_sprite[0][24][20] = 1; platform_sprite[0][24][21] = 1; platform_sprite[0][24][22] = 1; platform_sprite[0][24][23] = 1; platform_sprite[0][24][24] = 1; platform_sprite[0][25][5] = 1; platform_sprite[0][25][6] = 1; platform_sprite[0][25][7] = 1; platform_sprite[0][25][8] = 1; platform_sprite[0][25][9] = 1; platform_sprite[0][25][20] = 1; platform_sprite[0][25][21] = 1; platform_sprite[0][25][22] = 1; platform_sprite[0][25][23] = 1; platform_sprite[0][25][24] = 1; platform_sprite[0][26][5] = 1; platform_sprite[0][26][6] = 1; platform_sprite[0][26][7] = 1; platform_sprite[0][26][8] = 1; platform_sprite[0][26][9] = 1; platform_sprite[0][26][20] = 1; platform_sprite[0][26][21] = 1; platform_sprite[0][26][22] = 1; platform_sprite[0][26][23] = 1; platform_sprite[0][26][24] = 1; platform_sprite[0][27][5] = 1; platform_sprite[0][27][6] = 1; platform_sprite[0][27][7] = 1; platform_sprite[0][27][8] = 1; platform_sprite[0][27][9] = 1; platform_sprite[0][27][20] = 1; platform_sprite[0][27][21] = 1; platform_sprite[0][27][22] = 1; platform_sprite[0][27][23] = 1; platform_sprite[0][27][24] = 1; platform_sprite[0][28][5] = 1; platform_sprite[0][28][6] = 1; platform_sprite[0][28][7] = 1; platform_sprite[0][28][8] = 1; platform_sprite[0][28][9] = 1; platform_sprite[0][28][20] = 1; platform_sprite[0][28][21] = 1; platform_sprite[0][28][22] = 1; platform_sprite[0][28][23] = 1; platform_sprite[0][28][24] = 1; platform_sprite[0][29][5] = 1; platform_sprite[0][29][6] = 1; platform_sprite[0][29][7] = 1; platform_sprite[0][29][8] = 1; platform_sprite[0][29][9] = 1; platform_sprite[0][29][20] = 1; platform_sprite[0][29][21] = 1; platform_sprite[0][29][22] = 1; platform_sprite[0][29][23] = 1; platform_sprite[0][29][24] = 1; platform_sprite[0][30][5] = 1; platform_sprite[0][30][6] = 1; platform_sprite[0][30][7] = 1; platform_sprite[0][30][8] = 1; platform_sprite[0][30][9] = 1; platform_sprite[0][30][20] = 1; platform_sprite[0][30][21] = 1; platform_sprite[0][30][22] = 1; platform_sprite[0][30][23] = 1; platform_sprite[0][30][24] = 1; platform_sprite[0][31][5] = 1; platform_sprite[0][31][6] = 1; platform_sprite[0][31][7] = 1; platform_sprite[0][31][8] = 1; platform_sprite[0][31][9] = 1; platform_sprite[0][31][20] = 1; platform_sprite[0][31][21] = 1; platform_sprite[0][31][22] = 1; platform_sprite[0][31][23] = 1; platform_sprite[0][31][24] = 1; platform_sprite[0][32][5] = 1; platform_sprite[0][32][6] = 1; platform_sprite[0][32][7] = 1; platform_sprite[0][32][8] = 1; platform_sprite[0][32][9] = 1; platform_sprite[0][32][20] = 1; platform_sprite[0][32][21] = 1; platform_sprite[0][32][22] = 1; platform_sprite[0][32][23] = 1; platform_sprite[0][32][24] = 1; platform_sprite[0][33][5] = 1; platform_sprite[0][33][6] = 1; platform_sprite[0][33][7] = 1; platform_sprite[0][33][8] = 1; platform_sprite[0][33][9] = 1; platform_sprite[0][33][20] = 1; platform_sprite[0][33][21] = 1; platform_sprite[0][33][22] = 1; platform_sprite[0][33][23] = 1; platform_sprite[0][33][24] = 1; platform_sprite[0][34][5] = 1; platform_sprite[0][34][6] = 1; platform_sprite[0][34][7] = 1; platform_sprite[0][34][8] = 1; platform_sprite[0][34][9] = 1; platform_sprite[0][34][20] = 1; platform_sprite[0][34][21] = 1; platform_sprite[0][34][22] = 1; platform_sprite[0][34][23] = 1; platform_sprite[0][34][24] = 1; platform_sprite[0][35][5] = 1; platform_sprite[0][35][6] = 1; platform_sprite[0][35][7] = 1; platform_sprite[0][35][8] = 1; platform_sprite[0][35][9] = 1; platform_sprite[0][35][20] = 1; platform_sprite[0][35][21] = 1; platform_sprite[0][35][22] = 1; platform_sprite[0][35][23] = 1; platform_sprite[0][35][24] = 1; platform_sprite[0][36][5] = 1; platform_sprite[0][36][6] = 1; platform_sprite[0][36][7] = 1; platform_sprite[0][36][8] = 1; platform_sprite[0][36][9] = 1; platform_sprite[0][36][20] = 1; platform_sprite[0][36][21] = 1; platform_sprite[0][36][22] = 1; platform_sprite[0][36][23] = 1; platform_sprite[0][36][24] = 1; platform_sprite[0][37][5] = 1; platform_sprite[0][37][6] = 1; platform_sprite[0][37][7] = 1; platform_sprite[0][37][8] = 1; platform_sprite[0][37][9] = 1; platform_sprite[0][37][20] = 1; platform_sprite[0][37][21] = 1; platform_sprite[0][37][22] = 1; platform_sprite[0][37][23] = 1; platform_sprite[0][37][24] = 1; platform_sprite[0][38][5] = 1; platform_sprite[0][38][6] = 1; platform_sprite[0][38][7] = 1; platform_sprite[0][38][8] = 1; platform_sprite[0][38][9] = 1; platform_sprite[0][38][20] = 1; platform_sprite[0][38][21] = 1; platform_sprite[0][38][22] = 1; platform_sprite[0][38][23] = 1; platform_sprite[0][38][24] = 1; platform_sprite[0][39][5] = 1; platform_sprite[0][39][6] = 1; platform_sprite[0][39][7] = 1; platform_sprite[0][39][8] = 1; platform_sprite[0][39][9] = 1; platform_sprite[0][39][20] = 1; platform_sprite[0][39][21] = 1; platform_sprite[0][39][22] = 1; platform_sprite[0][39][23] = 1; platform_sprite[0][39][24] = 1; platform_sprite[0][40][5] = 1; platform_sprite[0][40][6] = 1; platform_sprite[0][40][7] = 1; platform_sprite[0][40][8] = 1; platform_sprite[0][40][9] = 1; platform_sprite[0][40][20] = 1; platform_sprite[0][40][21] = 1; platform_sprite[0][40][22] = 1; platform_sprite[0][40][23] = 1; platform_sprite[0][40][24] = 1; platform_sprite[0][41][5] = 1; platform_sprite[0][41][6] = 1; platform_sprite[0][41][7] = 1; platform_sprite[0][41][8] = 1; platform_sprite[0][41][9] = 1; platform_sprite[0][41][20] = 1; platform_sprite[0][41][21] = 1; platform_sprite[0][41][22] = 1; platform_sprite[0][41][23] = 1; platform_sprite[0][41][24] = 1; platform_sprite[0][42][5] = 1; platform_sprite[0][42][6] = 1; platform_sprite[0][42][7] = 1; platform_sprite[0][42][8] = 1; platform_sprite[0][42][9] = 1; platform_sprite[0][42][20] = 1; platform_sprite[0][42][21] = 1; platform_sprite[0][42][22] = 1; platform_sprite[0][42][23] = 1; platform_sprite[0][42][24] = 1; platform_sprite[0][43][5] = 1; platform_sprite[0][43][6] = 1; platform_sprite[0][43][7] = 1; platform_sprite[0][43][8] = 1; platform_sprite[0][43][9] = 1; platform_sprite[0][43][20] = 1; platform_sprite[0][43][21] = 1; platform_sprite[0][43][22] = 1; platform_sprite[0][43][23] = 1; platform_sprite[0][43][24] = 1; platform_sprite[0][44][5] = 1; platform_sprite[0][44][6] = 1; platform_sprite[0][44][7] = 1; platform_sprite[0][44][8] = 1; platform_sprite[0][44][9] = 1; platform_sprite[0][44][20] = 1; platform_sprite[0][44][21] = 1; platform_sprite[0][44][22] = 1; platform_sprite[0][44][23] = 1; platform_sprite[0][44][24] = 1; platform_sprite[0][45][5] = 1; platform_sprite[0][45][6] = 1; platform_sprite[0][45][7] = 1; platform_sprite[0][45][8] = 1; platform_sprite[0][45][9] = 1; platform_sprite[0][45][20] = 1; platform_sprite[0][45][21] = 1; platform_sprite[0][45][22] = 1; platform_sprite[0][45][23] = 1; platform_sprite[0][45][24] = 1; platform_sprite[0][46][5] = 1; platform_sprite[0][46][6] = 1; platform_sprite[0][46][7] = 1; platform_sprite[0][46][8] = 1; platform_sprite[0][46][9] = 1; platform_sprite[0][46][20] = 1; platform_sprite[0][46][21] = 1; platform_sprite[0][46][22] = 1; platform_sprite[0][46][23] = 1; platform_sprite[0][46][24] = 1; platform_sprite[0][47][5] = 1; platform_sprite[0][47][6] = 1; platform_sprite[0][47][7] = 1; platform_sprite[0][47][8] = 1; platform_sprite[0][47][9] = 1; platform_sprite[0][47][20] = 1; platform_sprite[0][47][21] = 1; platform_sprite[0][47][22] = 1; platform_sprite[0][47][23] = 1; platform_sprite[0][47][24] = 1; platform_sprite[0][48][5] = 1; platform_sprite[0][48][6] = 1; platform_sprite[0][48][7] = 1; platform_sprite[0][48][8] = 1; platform_sprite[0][48][9] = 1; platform_sprite[0][48][20] = 1; platform_sprite[0][48][21] = 1; platform_sprite[0][48][22] = 1; platform_sprite[0][48][23] = 1; platform_sprite[0][48][24] = 1; platform_sprite[0][49][5] = 1; platform_sprite[0][49][6] = 1; platform_sprite[0][49][7] = 1; platform_sprite[0][49][8] = 1; platform_sprite[0][49][9] = 1; platform_sprite[0][49][20] = 1; platform_sprite[0][49][21] = 1; platform_sprite[0][49][22] = 1; platform_sprite[0][49][23] = 1; platform_sprite[0][49][24] = 1; platform_sprite[0][50][5] = 1; platform_sprite[0][50][6] = 1; platform_sprite[0][50][7] = 1; platform_sprite[0][50][8] = 1; platform_sprite[0][50][9] = 1; platform_sprite[0][50][20] = 1; platform_sprite[0][50][21] = 1; platform_sprite[0][50][22] = 1; platform_sprite[0][50][23] = 1; platform_sprite[0][50][24] = 1; platform_sprite[0][51][5] = 1; platform_sprite[0][51][6] = 1; platform_sprite[0][51][7] = 1; platform_sprite[0][51][8] = 1; platform_sprite[0][51][9] = 1; platform_sprite[0][51][20] = 1; platform_sprite[0][51][21] = 1; platform_sprite[0][51][22] = 1; platform_sprite[0][51][23] = 1; platform_sprite[0][51][24] = 1; platform_sprite[0][52][5] = 1; platform_sprite[0][52][6] = 1; platform_sprite[0][52][7] = 1; platform_sprite[0][52][8] = 1; platform_sprite[0][52][9] = 1; platform_sprite[0][52][20] = 1; platform_sprite[0][52][21] = 1; platform_sprite[0][52][22] = 1; platform_sprite[0][52][23] = 1; platform_sprite[0][52][24] = 1; platform_sprite[0][53][5] = 1; platform_sprite[0][53][6] = 1; platform_sprite[0][53][7] = 1; platform_sprite[0][53][8] = 1; platform_sprite[0][53][9] = 1; platform_sprite[0][53][20] = 1; platform_sprite[0][53][21] = 1; platform_sprite[0][53][22] = 1; platform_sprite[0][53][23] = 1; platform_sprite[0][53][24] = 1; platform_sprite[0][54][5] = 1; platform_sprite[0][54][6] = 1; platform_sprite[0][54][7] = 1; platform_sprite[0][54][8] = 1; platform_sprite[0][54][9] = 1; platform_sprite[0][54][20] = 1; platform_sprite[0][54][21] = 1; platform_sprite[0][54][22] = 1; platform_sprite[0][54][23] = 1; platform_sprite[0][54][24] = 1; platform_sprite[0][55][5] = 1; platform_sprite[0][55][6] = 1; platform_sprite[0][55][7] = 1; platform_sprite[0][55][8] = 1; platform_sprite[0][55][9] = 1; platform_sprite[0][55][20] = 1; platform_sprite[0][55][21] = 1; platform_sprite[0][55][22] = 1; platform_sprite[0][55][23] = 1; platform_sprite[0][55][24] = 1; platform_sprite[0][56][5] = 1; platform_sprite[0][56][6] = 1; platform_sprite[0][56][7] = 1; platform_sprite[0][56][8] = 1; platform_sprite[0][56][9] = 1; platform_sprite[0][56][20] = 1; platform_sprite[0][56][21] = 1; platform_sprite[0][56][22] = 1; platform_sprite[0][56][23] = 1; platform_sprite[0][56][24] = 1; platform_sprite[0][57][5] = 1; platform_sprite[0][57][6] = 1; platform_sprite[0][57][7] = 1; platform_sprite[0][57][8] = 1; platform_sprite[0][57][9] = 1; platform_sprite[0][57][20] = 1; platform_sprite[0][57][21] = 1; platform_sprite[0][57][22] = 1; platform_sprite[0][57][23] = 1; platform_sprite[0][57][24] = 1; platform_sprite[0][58][5] = 1; platform_sprite[0][58][6] = 1; platform_sprite[0][58][7] = 1; platform_sprite[0][58][8] = 1; platform_sprite[0][58][9] = 1; platform_sprite[0][58][20] = 1; platform_sprite[0][58][21] = 1; platform_sprite[0][58][22] = 1; platform_sprite[0][58][23] = 1; platform_sprite[0][58][24] = 1; platform_sprite[0][59][5] = 1; platform_sprite[0][59][6] = 1; platform_sprite[0][59][7] = 1; platform_sprite[0][59][8] = 1; platform_sprite[0][59][9] = 1; platform_sprite[0][59][20] = 1; platform_sprite[0][59][21] = 1; platform_sprite[0][59][22] = 1; platform_sprite[0][59][23] = 1; platform_sprite[0][59][24] = 1; platform_sprite[0][60][5] = 1; platform_sprite[0][60][6] = 1; platform_sprite[0][60][7] = 1; platform_sprite[0][60][8] = 1; platform_sprite[0][60][9] = 1; platform_sprite[0][60][20] = 1; platform_sprite[0][60][21] = 1; platform_sprite[0][60][22] = 1; platform_sprite[0][60][23] = 1; platform_sprite[0][60][24] = 1; platform_sprite[0][61][5] = 1; platform_sprite[0][61][6] = 1; platform_sprite[0][61][7] = 1; platform_sprite[0][61][8] = 1; platform_sprite[0][61][9] = 1; platform_sprite[0][61][20] = 1; platform_sprite[0][61][21] = 1; platform_sprite[0][61][22] = 1; platform_sprite[0][61][23] = 1; platform_sprite[0][61][24] = 1; platform_sprite[0][62][5] = 1; platform_sprite[0][62][6] = 1; platform_sprite[0][62][7] = 1; platform_sprite[0][62][8] = 1; platform_sprite[0][62][9] = 1; platform_sprite[0][62][20] = 1; platform_sprite[0][62][21] = 1; platform_sprite[0][62][22] = 1; platform_sprite[0][62][23] = 1; platform_sprite[0][62][24] = 1; platform_sprite[0][63][5] = 1; platform_sprite[0][63][6] = 1; platform_sprite[0][63][7] = 1; platform_sprite[0][63][8] = 1; platform_sprite[0][63][9] = 1; platform_sprite[0][63][20] = 1; platform_sprite[0][63][21] = 1; platform_sprite[0][63][22] = 1; platform_sprite[0][63][23] = 1; platform_sprite[0][63][24] = 1; platform_sprite[0][64][5] = 1; platform_sprite[0][64][6] = 1; platform_sprite[0][64][7] = 1; platform_sprite[0][64][8] = 1; platform_sprite[0][64][9] = 1; platform_sprite[0][64][20] = 1; platform_sprite[0][64][21] = 1; platform_sprite[0][64][22] = 1; platform_sprite[0][64][23] = 1; platform_sprite[0][64][24] = 1; platform_sprite[0][65][5] = 1; platform_sprite[0][65][6] = 1; platform_sprite[0][65][7] = 1; platform_sprite[0][65][8] = 1; platform_sprite[0][65][9] = 1; platform_sprite[0][65][20] = 1; platform_sprite[0][65][21] = 1; platform_sprite[0][65][22] = 1; platform_sprite[0][65][23] = 1; platform_sprite[0][65][24] = 1; platform_sprite[0][66][5] = 1; platform_sprite[0][66][6] = 1; platform_sprite[0][66][7] = 1; platform_sprite[0][66][8] = 1; platform_sprite[0][66][9] = 1; platform_sprite[0][66][20] = 1; platform_sprite[0][66][21] = 1; platform_sprite[0][66][22] = 1; platform_sprite[0][66][23] = 1; platform_sprite[0][66][24] = 1; platform_sprite[0][67][5] = 1; platform_sprite[0][67][6] = 1; platform_sprite[0][67][7] = 1; platform_sprite[0][67][8] = 1; platform_sprite[0][67][9] = 1; platform_sprite[0][67][20] = 1; platform_sprite[0][67][21] = 1; platform_sprite[0][67][22] = 1; platform_sprite[0][67][23] = 1; platform_sprite[0][67][24] = 1; platform_sprite[0][68][5] = 1; platform_sprite[0][68][6] = 1; platform_sprite[0][68][7] = 1; platform_sprite[0][68][8] = 1; platform_sprite[0][68][9] = 1; platform_sprite[0][68][20] = 1; platform_sprite[0][68][21] = 1; platform_sprite[0][68][22] = 1; platform_sprite[0][68][23] = 1; platform_sprite[0][68][24] = 1; platform_sprite[0][69][5] = 1; platform_sprite[0][69][6] = 1; platform_sprite[0][69][7] = 1; platform_sprite[0][69][8] = 1; platform_sprite[0][69][9] = 1; platform_sprite[0][69][20] = 1; platform_sprite[0][69][21] = 1; platform_sprite[0][69][22] = 1; platform_sprite[0][69][23] = 1; platform_sprite[0][69][24] = 1; platform_sprite[0][70][5] = 1; platform_sprite[0][70][6] = 1; platform_sprite[0][70][7] = 1; platform_sprite[0][70][8] = 1; platform_sprite[0][70][9] = 1; platform_sprite[0][70][20] = 1; platform_sprite[0][70][21] = 1; platform_sprite[0][70][22] = 1; platform_sprite[0][70][23] = 1; platform_sprite[0][70][24] = 1; platform_sprite[0][71][5] = 1; platform_sprite[0][71][6] = 1; platform_sprite[0][71][7] = 1; platform_sprite[0][71][8] = 1; platform_sprite[0][71][9] = 1; platform_sprite[0][71][20] = 1; platform_sprite[0][71][21] = 1; platform_sprite[0][71][22] = 1; platform_sprite[0][71][23] = 1; platform_sprite[0][71][24] = 1; platform_sprite[0][72][5] = 1; platform_sprite[0][72][6] = 1; platform_sprite[0][72][7] = 1; platform_sprite[0][72][8] = 1; platform_sprite[0][72][9] = 1; platform_sprite[0][72][20] = 1; platform_sprite[0][72][21] = 1; platform_sprite[0][72][22] = 1; platform_sprite[0][72][23] = 1; platform_sprite[0][72][24] = 1; platform_sprite[0][73][5] = 1; platform_sprite[0][73][6] = 1; platform_sprite[0][73][7] = 1; platform_sprite[0][73][8] = 1; platform_sprite[0][73][9] = 1; platform_sprite[0][73][20] = 1; platform_sprite[0][73][21] = 1; platform_sprite[0][73][22] = 1; platform_sprite[0][73][23] = 1; platform_sprite[0][73][24] = 1; platform_sprite[0][74][5] = 1; platform_sprite[0][74][6] = 1; platform_sprite[0][74][7] = 1; platform_sprite[0][74][8] = 1; platform_sprite[0][74][9] = 1; platform_sprite[0][74][20] = 1; platform_sprite[0][74][21] = 1; platform_sprite[0][74][22] = 1; platform_sprite[0][74][23] = 1; platform_sprite[0][74][24] = 1; platform_sprite[0][75][5] = 1; platform_sprite[0][75][6] = 1; platform_sprite[0][75][7] = 1; platform_sprite[0][75][8] = 1; platform_sprite[0][75][9] = 1; platform_sprite[0][75][20] = 1; platform_sprite[0][75][21] = 1; platform_sprite[0][75][22] = 1; platform_sprite[0][75][23] = 1; platform_sprite[0][75][24] = 1; platform_sprite[0][76][5] = 1; platform_sprite[0][76][6] = 1; platform_sprite[0][76][7] = 1; platform_sprite[0][76][8] = 1; platform_sprite[0][76][9] = 1; platform_sprite[0][76][20] = 1; platform_sprite[0][76][21] = 1; platform_sprite[0][76][22] = 1; platform_sprite[0][76][23] = 1; platform_sprite[0][76][24] = 1; platform_sprite[0][77][5] = 1; platform_sprite[0][77][6] = 1; platform_sprite[0][77][7] = 1; platform_sprite[0][77][8] = 1; platform_sprite[0][77][9] = 1; platform_sprite[0][77][20] = 1; platform_sprite[0][77][21] = 1; platform_sprite[0][77][22] = 1; platform_sprite[0][77][23] = 1; platform_sprite[0][77][24] = 1; platform_sprite[0][78][5] = 1; platform_sprite[0][78][6] = 1; platform_sprite[0][78][7] = 1; platform_sprite[0][78][8] = 1; platform_sprite[0][78][9] = 1; platform_sprite[0][78][20] = 1; platform_sprite[0][78][21] = 1; platform_sprite[0][78][22] = 1; platform_sprite[0][78][23] = 1; platform_sprite[0][78][24] = 1; platform_sprite[0][79][5] = 1; platform_sprite[0][79][6] = 1; platform_sprite[0][79][7] = 1; platform_sprite[0][79][8] = 1; platform_sprite[0][79][9] = 1; platform_sprite[0][79][20] = 1; platform_sprite[0][79][21] = 1; platform_sprite[0][79][22] = 1; platform_sprite[0][79][23] = 1; platform_sprite[0][79][24] = 1; platform_sprite[0][80][5] = 1; platform_sprite[0][80][6] = 1; platform_sprite[0][80][7] = 1; platform_sprite[0][80][8] = 1; platform_sprite[0][80][9] = 1; platform_sprite[0][80][20] = 1; platform_sprite[0][80][21] = 1; platform_sprite[0][80][22] = 1; platform_sprite[0][80][23] = 1; platform_sprite[0][80][24] = 1; platform_sprite[0][81][5] = 1; platform_sprite[0][81][6] = 1; platform_sprite[0][81][7] = 1; platform_sprite[0][81][8] = 1; platform_sprite[0][81][9] = 1; platform_sprite[0][81][20] = 1; platform_sprite[0][81][21] = 1; platform_sprite[0][81][22] = 1; platform_sprite[0][81][23] = 1; platform_sprite[0][81][24] = 1; platform_sprite[0][82][5] = 1; platform_sprite[0][82][6] = 1; platform_sprite[0][82][7] = 1; platform_sprite[0][82][8] = 1; platform_sprite[0][82][9] = 1; platform_sprite[0][82][20] = 1; platform_sprite[0][82][21] = 1; platform_sprite[0][82][22] = 1; platform_sprite[0][82][23] = 1; platform_sprite[0][82][24] = 1; platform_sprite[0][83][5] = 1; platform_sprite[0][83][6] = 1; platform_sprite[0][83][7] = 1; platform_sprite[0][83][8] = 1; platform_sprite[0][83][9] = 1; platform_sprite[0][83][20] = 1; platform_sprite[0][83][21] = 1; platform_sprite[0][83][22] = 1; platform_sprite[0][83][23] = 1; platform_sprite[0][83][24] = 1; platform_sprite[0][84][5] = 1; platform_sprite[0][84][6] = 1; platform_sprite[0][84][7] = 1; platform_sprite[0][84][8] = 1; platform_sprite[0][84][9] = 1; platform_sprite[0][84][20] = 1; platform_sprite[0][84][21] = 1; platform_sprite[0][84][22] = 1; platform_sprite[0][84][23] = 1; platform_sprite[0][84][24] = 1; platform_sprite[0][85][5] = 1; platform_sprite[0][85][6] = 1; platform_sprite[0][85][7] = 1; platform_sprite[0][85][8] = 1; platform_sprite[0][85][9] = 1; platform_sprite[0][85][20] = 1; platform_sprite[0][85][21] = 1; platform_sprite[0][85][22] = 1; platform_sprite[0][85][23] = 1; platform_sprite[0][85][24] = 1; platform_sprite[0][86][5] = 1; platform_sprite[0][86][6] = 1; platform_sprite[0][86][7] = 1; platform_sprite[0][86][8] = 1; platform_sprite[0][86][9] = 1; platform_sprite[0][86][20] = 1; platform_sprite[0][86][21] = 1; platform_sprite[0][86][22] = 1; platform_sprite[0][86][23] = 1; platform_sprite[0][86][24] = 1; platform_sprite[0][87][5] = 1; platform_sprite[0][87][6] = 1; platform_sprite[0][87][7] = 1; platform_sprite[0][87][8] = 1; platform_sprite[0][87][9] = 1; platform_sprite[0][87][20] = 1; platform_sprite[0][87][21] = 1; platform_sprite[0][87][22] = 1; platform_sprite[0][87][23] = 1; platform_sprite[0][87][24] = 1; platform_sprite[0][88][5] = 1; platform_sprite[0][88][6] = 1; platform_sprite[0][88][7] = 1; platform_sprite[0][88][8] = 1; platform_sprite[0][88][9] = 1; platform_sprite[0][88][20] = 1; platform_sprite[0][88][21] = 1; platform_sprite[0][88][22] = 1; platform_sprite[0][88][23] = 1; platform_sprite[0][88][24] = 1; platform_sprite[0][89][5] = 1; platform_sprite[0][89][6] = 1; platform_sprite[0][89][7] = 1; platform_sprite[0][89][8] = 1; platform_sprite[0][89][9] = 1; platform_sprite[0][89][20] = 1; platform_sprite[0][89][21] = 1; platform_sprite[0][89][22] = 1; platform_sprite[0][89][23] = 1; platform_sprite[0][89][24] = 1; platform_sprite[0][90][10] = 1; platform_sprite[0][90][11] = 1; platform_sprite[0][90][12] = 1; platform_sprite[0][90][13] = 1; platform_sprite[0][90][14] = 1; platform_sprite[0][90][15] = 1; platform_sprite[0][90][16] = 1; platform_sprite[0][90][17] = 1; platform_sprite[0][90][18] = 1; platform_sprite[0][90][19] = 1; platform_sprite[0][91][10] = 1; platform_sprite[0][91][11] = 1; platform_sprite[0][91][12] = 1; platform_sprite[0][91][13] = 1; platform_sprite[0][91][14] = 1; platform_sprite[0][91][15] = 1; platform_sprite[0][91][16] = 1; platform_sprite[0][91][17] = 1; platform_sprite[0][91][18] = 1; platform_sprite[0][91][19] = 1; platform_sprite[0][92][10] = 1; platform_sprite[0][92][11] = 1; platform_sprite[0][92][12] = 1; platform_sprite[0][92][13] = 1; platform_sprite[0][92][14] = 1; platform_sprite[0][92][15] = 1; platform_sprite[0][92][16] = 1; platform_sprite[0][92][17] = 1; platform_sprite[0][92][18] = 1; platform_sprite[0][92][19] = 1; platform_sprite[0][93][10] = 1; platform_sprite[0][93][11] = 1; platform_sprite[0][93][12] = 1; platform_sprite[0][93][13] = 1; platform_sprite[0][93][14] = 1; platform_sprite[0][93][15] = 1; platform_sprite[0][93][16] = 1; platform_sprite[0][93][17] = 1; platform_sprite[0][93][18] = 1; platform_sprite[0][93][19] = 1; platform_sprite[0][94][10] = 1; platform_sprite[0][94][11] = 1; platform_sprite[0][94][12] = 1; platform_sprite[0][94][13] = 1; platform_sprite[0][94][14] = 1; platform_sprite[0][94][15] = 1; platform_sprite[0][94][16] = 1; platform_sprite[0][94][17] = 1; platform_sprite[0][94][18] = 1; platform_sprite[0][94][19] = 1; 
					platform_sprite[1][5][10] = 1; platform_sprite[1][5][11] = 1; platform_sprite[1][5][12] = 1; platform_sprite[1][5][13] = 1; platform_sprite[1][5][14] = 1; platform_sprite[1][5][15] = 1; platform_sprite[1][5][16] = 1; platform_sprite[1][5][17] = 1; platform_sprite[1][5][18] = 1; platform_sprite[1][5][19] = 1; platform_sprite[1][6][10] = 1; platform_sprite[1][6][11] = 1; platform_sprite[1][6][12] = 1; platform_sprite[1][6][13] = 1; platform_sprite[1][6][14] = 1; platform_sprite[1][6][15] = 1; platform_sprite[1][6][16] = 1; platform_sprite[1][6][17] = 1; platform_sprite[1][6][18] = 1; platform_sprite[1][6][19] = 1; platform_sprite[1][7][10] = 1; platform_sprite[1][7][11] = 1; platform_sprite[1][7][12] = 1; platform_sprite[1][7][13] = 1; platform_sprite[1][7][14] = 1; platform_sprite[1][7][15] = 1; platform_sprite[1][7][16] = 1; platform_sprite[1][7][17] = 1; platform_sprite[1][7][18] = 1; platform_sprite[1][7][19] = 1; platform_sprite[1][8][10] = 1; platform_sprite[1][8][11] = 1; platform_sprite[1][8][12] = 1; platform_sprite[1][8][13] = 1; platform_sprite[1][8][14] = 1; platform_sprite[1][8][15] = 1; platform_sprite[1][8][16] = 1; platform_sprite[1][8][17] = 1; platform_sprite[1][8][18] = 1; platform_sprite[1][8][19] = 1; platform_sprite[1][9][10] = 1; platform_sprite[1][9][11] = 1; platform_sprite[1][9][12] = 1; platform_sprite[1][9][13] = 1; platform_sprite[1][9][14] = 1; platform_sprite[1][9][15] = 1; platform_sprite[1][9][16] = 1; platform_sprite[1][9][17] = 1; platform_sprite[1][9][18] = 1; platform_sprite[1][9][19] = 1; platform_sprite[1][9][20] = 1; platform_sprite[1][9][21] = 1; platform_sprite[1][9][22] = 1; platform_sprite[1][9][23] = 1; platform_sprite[1][9][24] = 1; platform_sprite[1][10][5] = 1; platform_sprite[1][10][6] = 1; platform_sprite[1][10][7] = 1; platform_sprite[1][10][8] = 1; platform_sprite[1][10][9] = 1; platform_sprite[1][10][20] = 1; platform_sprite[1][10][21] = 1; platform_sprite[1][10][22] = 1; platform_sprite[1][10][23] = 1; platform_sprite[1][10][24] = 1; platform_sprite[1][11][5] = 1; platform_sprite[1][11][6] = 1; platform_sprite[1][11][7] = 1; platform_sprite[1][11][8] = 1; platform_sprite[1][11][9] = 1; platform_sprite[1][11][20] = 1; platform_sprite[1][11][21] = 1; platform_sprite[1][11][22] = 1; platform_sprite[1][11][23] = 1; platform_sprite[1][11][24] = 1; platform_sprite[1][12][5] = 1; platform_sprite[1][12][6] = 1; platform_sprite[1][12][7] = 1; platform_sprite[1][12][8] = 1; platform_sprite[1][12][9] = 1; platform_sprite[1][12][20] = 1; platform_sprite[1][12][21] = 1; platform_sprite[1][12][22] = 1; platform_sprite[1][12][23] = 1; platform_sprite[1][12][24] = 1; platform_sprite[1][13][5] = 1; platform_sprite[1][13][6] = 1; platform_sprite[1][13][7] = 1; platform_sprite[1][13][8] = 1; platform_sprite[1][13][9] = 1; platform_sprite[1][13][20] = 1; platform_sprite[1][13][21] = 1; platform_sprite[1][13][22] = 1; platform_sprite[1][13][23] = 1; platform_sprite[1][13][24] = 1; platform_sprite[1][14][5] = 1; platform_sprite[1][14][6] = 1; platform_sprite[1][14][7] = 1; platform_sprite[1][14][8] = 1; platform_sprite[1][14][9] = 1; platform_sprite[1][14][20] = 1; platform_sprite[1][14][21] = 1; platform_sprite[1][14][22] = 1; platform_sprite[1][14][23] = 1; platform_sprite[1][14][24] = 1; platform_sprite[1][15][5] = 1; platform_sprite[1][15][6] = 1; platform_sprite[1][15][7] = 1; platform_sprite[1][15][8] = 1; platform_sprite[1][15][9] = 1; platform_sprite[1][15][20] = 1; platform_sprite[1][15][21] = 1; platform_sprite[1][15][22] = 1; platform_sprite[1][15][23] = 1; platform_sprite[1][15][24] = 1; platform_sprite[1][16][5] = 1; platform_sprite[1][16][6] = 1; platform_sprite[1][16][7] = 1; platform_sprite[1][16][8] = 1; platform_sprite[1][16][9] = 1; platform_sprite[1][16][20] = 1; platform_sprite[1][16][21] = 1; platform_sprite[1][16][22] = 1; platform_sprite[1][16][23] = 1; platform_sprite[1][16][24] = 1; platform_sprite[1][17][5] = 1; platform_sprite[1][17][6] = 1; platform_sprite[1][17][7] = 1; platform_sprite[1][17][8] = 1; platform_sprite[1][17][9] = 1; platform_sprite[1][17][20] = 1; platform_sprite[1][17][21] = 1; platform_sprite[1][17][22] = 1; platform_sprite[1][17][23] = 1; platform_sprite[1][17][24] = 1; platform_sprite[1][18][5] = 1; platform_sprite[1][18][6] = 1; platform_sprite[1][18][7] = 1; platform_sprite[1][18][8] = 1; platform_sprite[1][18][9] = 1; platform_sprite[1][18][20] = 1; platform_sprite[1][18][21] = 1; platform_sprite[1][18][22] = 1; platform_sprite[1][18][23] = 1; platform_sprite[1][18][24] = 1; platform_sprite[1][19][5] = 1; platform_sprite[1][19][6] = 1; platform_sprite[1][19][7] = 1; platform_sprite[1][19][8] = 1; platform_sprite[1][19][9] = 1; platform_sprite[1][19][20] = 1; platform_sprite[1][19][21] = 1; platform_sprite[1][19][22] = 1; platform_sprite[1][19][23] = 1; platform_sprite[1][19][24] = 1; platform_sprite[1][20][5] = 1; platform_sprite[1][20][6] = 1; platform_sprite[1][20][7] = 1; platform_sprite[1][20][8] = 1; platform_sprite[1][20][9] = 1; platform_sprite[1][20][20] = 1; platform_sprite[1][20][21] = 1; platform_sprite[1][20][22] = 1; platform_sprite[1][20][23] = 1; platform_sprite[1][20][24] = 1; platform_sprite[1][21][5] = 1; platform_sprite[1][21][6] = 1; platform_sprite[1][21][7] = 1; platform_sprite[1][21][8] = 1; platform_sprite[1][21][9] = 1; platform_sprite[1][21][20] = 1; platform_sprite[1][21][21] = 1; platform_sprite[1][21][22] = 1; platform_sprite[1][21][23] = 1; platform_sprite[1][21][24] = 1; platform_sprite[1][22][5] = 1; platform_sprite[1][22][6] = 1; platform_sprite[1][22][7] = 1; platform_sprite[1][22][8] = 1; platform_sprite[1][22][9] = 1; platform_sprite[1][22][20] = 1; platform_sprite[1][22][21] = 1; platform_sprite[1][22][22] = 1; platform_sprite[1][22][23] = 1; platform_sprite[1][22][24] = 1; platform_sprite[1][23][5] = 1; platform_sprite[1][23][6] = 1; platform_sprite[1][23][7] = 1; platform_sprite[1][23][8] = 1; platform_sprite[1][23][9] = 1; platform_sprite[1][23][20] = 1; platform_sprite[1][23][21] = 1; platform_sprite[1][23][22] = 1; platform_sprite[1][23][23] = 1; platform_sprite[1][23][24] = 1; platform_sprite[1][24][5] = 1; platform_sprite[1][24][6] = 1; platform_sprite[1][24][7] = 1; platform_sprite[1][24][8] = 1; platform_sprite[1][24][9] = 1; platform_sprite[1][24][20] = 1; platform_sprite[1][24][21] = 1; platform_sprite[1][24][22] = 1; platform_sprite[1][24][23] = 1; platform_sprite[1][24][24] = 1; platform_sprite[1][25][5] = 1; platform_sprite[1][25][6] = 1; platform_sprite[1][25][7] = 1; platform_sprite[1][25][8] = 1; platform_sprite[1][25][9] = 1; platform_sprite[1][25][20] = 1; platform_sprite[1][25][21] = 1; platform_sprite[1][25][22] = 1; platform_sprite[1][25][23] = 1; platform_sprite[1][25][24] = 1; platform_sprite[1][26][5] = 1; platform_sprite[1][26][6] = 1; platform_sprite[1][26][7] = 1; platform_sprite[1][26][8] = 1; platform_sprite[1][26][9] = 1; platform_sprite[1][26][20] = 1; platform_sprite[1][26][21] = 1; platform_sprite[1][26][22] = 1; platform_sprite[1][26][23] = 1; platform_sprite[1][26][24] = 1; platform_sprite[1][27][5] = 1; platform_sprite[1][27][6] = 1; platform_sprite[1][27][7] = 1; platform_sprite[1][27][8] = 1; platform_sprite[1][27][9] = 1; platform_sprite[1][27][20] = 1; platform_sprite[1][27][21] = 1; platform_sprite[1][27][22] = 1; platform_sprite[1][27][23] = 1; platform_sprite[1][27][24] = 1; platform_sprite[1][28][5] = 1; platform_sprite[1][28][6] = 1; platform_sprite[1][28][7] = 1; platform_sprite[1][28][8] = 1; platform_sprite[1][28][9] = 1; platform_sprite[1][28][20] = 1; platform_sprite[1][28][21] = 1; platform_sprite[1][28][22] = 1; platform_sprite[1][28][23] = 1; platform_sprite[1][28][24] = 1; platform_sprite[1][29][5] = 1; platform_sprite[1][29][6] = 1; platform_sprite[1][29][7] = 1; platform_sprite[1][29][8] = 1; platform_sprite[1][29][9] = 1; platform_sprite[1][29][20] = 1; platform_sprite[1][29][21] = 1; platform_sprite[1][29][22] = 1; platform_sprite[1][29][23] = 1; platform_sprite[1][29][24] = 1; platform_sprite[1][30][5] = 1; platform_sprite[1][30][6] = 1; platform_sprite[1][30][7] = 1; platform_sprite[1][30][8] = 1; platform_sprite[1][30][9] = 1; platform_sprite[1][30][20] = 1; platform_sprite[1][30][21] = 1; platform_sprite[1][30][22] = 1; platform_sprite[1][30][23] = 1; platform_sprite[1][30][24] = 1; platform_sprite[1][31][5] = 1; platform_sprite[1][31][6] = 1; platform_sprite[1][31][7] = 1; platform_sprite[1][31][8] = 1; platform_sprite[1][31][9] = 1; platform_sprite[1][31][20] = 1; platform_sprite[1][31][21] = 1; platform_sprite[1][31][22] = 1; platform_sprite[1][31][23] = 1; platform_sprite[1][31][24] = 1; platform_sprite[1][32][5] = 1; platform_sprite[1][32][6] = 1; platform_sprite[1][32][7] = 1; platform_sprite[1][32][8] = 1; platform_sprite[1][32][9] = 1; platform_sprite[1][32][20] = 1; platform_sprite[1][32][21] = 1; platform_sprite[1][32][22] = 1; platform_sprite[1][32][23] = 1; platform_sprite[1][32][24] = 1; platform_sprite[1][33][5] = 1; platform_sprite[1][33][6] = 1; platform_sprite[1][33][7] = 1; platform_sprite[1][33][8] = 1; platform_sprite[1][33][9] = 1; platform_sprite[1][33][20] = 1; platform_sprite[1][33][21] = 1; platform_sprite[1][33][22] = 1; platform_sprite[1][33][23] = 1; platform_sprite[1][33][24] = 1; platform_sprite[1][34][5] = 1; platform_sprite[1][34][6] = 1; platform_sprite[1][34][7] = 1; platform_sprite[1][34][8] = 1; platform_sprite[1][34][9] = 1; platform_sprite[1][34][20] = 1; platform_sprite[1][34][21] = 1; platform_sprite[1][34][22] = 1; platform_sprite[1][34][23] = 1; platform_sprite[1][34][24] = 1; platform_sprite[1][35][5] = 1; platform_sprite[1][35][6] = 1; platform_sprite[1][35][7] = 1; platform_sprite[1][35][8] = 1; platform_sprite[1][35][9] = 1; platform_sprite[1][35][20] = 1; platform_sprite[1][35][21] = 1; platform_sprite[1][35][22] = 1; platform_sprite[1][35][23] = 1; platform_sprite[1][35][24] = 1; platform_sprite[1][36][5] = 1; platform_sprite[1][36][6] = 1; platform_sprite[1][36][7] = 1; platform_sprite[1][36][8] = 1; platform_sprite[1][36][9] = 1; platform_sprite[1][36][20] = 1; platform_sprite[1][36][21] = 1; platform_sprite[1][36][22] = 1; platform_sprite[1][36][23] = 1; platform_sprite[1][36][24] = 1; platform_sprite[1][37][5] = 1; platform_sprite[1][37][6] = 1; platform_sprite[1][37][7] = 1; platform_sprite[1][37][8] = 1; platform_sprite[1][37][9] = 1; platform_sprite[1][37][20] = 1; platform_sprite[1][37][21] = 1; platform_sprite[1][37][22] = 1; platform_sprite[1][37][23] = 1; platform_sprite[1][37][24] = 1; platform_sprite[1][38][5] = 1; platform_sprite[1][38][6] = 1; platform_sprite[1][38][7] = 1; platform_sprite[1][38][8] = 1; platform_sprite[1][38][9] = 1; platform_sprite[1][38][20] = 1; platform_sprite[1][38][21] = 1; platform_sprite[1][38][22] = 1; platform_sprite[1][38][23] = 1; platform_sprite[1][38][24] = 1; platform_sprite[1][39][5] = 1; platform_sprite[1][39][6] = 1; platform_sprite[1][39][7] = 1; platform_sprite[1][39][8] = 1; platform_sprite[1][39][9] = 1; platform_sprite[1][39][20] = 1; platform_sprite[1][39][21] = 1; platform_sprite[1][39][22] = 1; platform_sprite[1][39][23] = 1; platform_sprite[1][39][24] = 1; platform_sprite[1][40][5] = 1; platform_sprite[1][40][6] = 1; platform_sprite[1][40][7] = 1; platform_sprite[1][40][8] = 1; platform_sprite[1][40][9] = 1; platform_sprite[1][40][20] = 1; platform_sprite[1][40][21] = 1; platform_sprite[1][40][22] = 1; platform_sprite[1][40][23] = 1; platform_sprite[1][40][24] = 1; platform_sprite[1][41][5] = 1; platform_sprite[1][41][6] = 1; platform_sprite[1][41][7] = 1; platform_sprite[1][41][8] = 1; platform_sprite[1][41][9] = 1; platform_sprite[1][41][20] = 1; platform_sprite[1][41][21] = 1; platform_sprite[1][41][22] = 1; platform_sprite[1][41][23] = 1; platform_sprite[1][41][24] = 1; platform_sprite[1][42][5] = 1; platform_sprite[1][42][6] = 1; platform_sprite[1][42][7] = 1; platform_sprite[1][42][8] = 1; platform_sprite[1][42][9] = 1; platform_sprite[1][42][20] = 1; platform_sprite[1][42][21] = 1; platform_sprite[1][42][22] = 1; platform_sprite[1][42][23] = 1; platform_sprite[1][42][24] = 1; platform_sprite[1][43][5] = 1; platform_sprite[1][43][6] = 1; platform_sprite[1][43][7] = 1; platform_sprite[1][43][8] = 1; platform_sprite[1][43][9] = 1; platform_sprite[1][43][20] = 1; platform_sprite[1][43][21] = 1; platform_sprite[1][43][22] = 1; platform_sprite[1][43][23] = 1; platform_sprite[1][43][24] = 1; platform_sprite[1][44][5] = 1; platform_sprite[1][44][6] = 1; platform_sprite[1][44][7] = 1; platform_sprite[1][44][8] = 1; platform_sprite[1][44][9] = 1; platform_sprite[1][44][20] = 1; platform_sprite[1][44][21] = 1; platform_sprite[1][44][22] = 1; platform_sprite[1][44][23] = 1; platform_sprite[1][44][24] = 1; platform_sprite[1][45][5] = 1; platform_sprite[1][45][6] = 1; platform_sprite[1][45][7] = 1; platform_sprite[1][45][8] = 1; platform_sprite[1][45][9] = 1; platform_sprite[1][45][20] = 1; platform_sprite[1][45][21] = 1; platform_sprite[1][45][22] = 1; platform_sprite[1][45][23] = 1; platform_sprite[1][45][24] = 1; platform_sprite[1][46][5] = 1; platform_sprite[1][46][6] = 1; platform_sprite[1][46][7] = 1; platform_sprite[1][46][8] = 1; platform_sprite[1][46][9] = 1; platform_sprite[1][46][20] = 1; platform_sprite[1][46][21] = 1; platform_sprite[1][46][22] = 1; platform_sprite[1][46][23] = 1; platform_sprite[1][46][24] = 1; platform_sprite[1][47][5] = 1; platform_sprite[1][47][6] = 1; platform_sprite[1][47][7] = 1; platform_sprite[1][47][8] = 1; platform_sprite[1][47][9] = 1; platform_sprite[1][47][20] = 1; platform_sprite[1][47][21] = 1; platform_sprite[1][47][22] = 1; platform_sprite[1][47][23] = 1; platform_sprite[1][47][24] = 1; platform_sprite[1][48][5] = 1; platform_sprite[1][48][6] = 1; platform_sprite[1][48][7] = 1; platform_sprite[1][48][8] = 1; platform_sprite[1][48][9] = 1; platform_sprite[1][48][20] = 1; platform_sprite[1][48][21] = 1; platform_sprite[1][48][22] = 1; platform_sprite[1][48][23] = 1; platform_sprite[1][48][24] = 1; platform_sprite[1][49][5] = 1; platform_sprite[1][49][6] = 1; platform_sprite[1][49][7] = 1; platform_sprite[1][49][8] = 1; platform_sprite[1][49][9] = 1; platform_sprite[1][49][20] = 1; platform_sprite[1][49][21] = 1; platform_sprite[1][49][22] = 1; platform_sprite[1][49][23] = 1; platform_sprite[1][49][24] = 1; platform_sprite[1][50][5] = 1; platform_sprite[1][50][6] = 1; platform_sprite[1][50][7] = 1; platform_sprite[1][50][8] = 1; platform_sprite[1][50][9] = 1; platform_sprite[1][50][20] = 1; platform_sprite[1][50][21] = 1; platform_sprite[1][50][22] = 1; platform_sprite[1][50][23] = 1; platform_sprite[1][50][24] = 1; platform_sprite[1][51][5] = 1; platform_sprite[1][51][6] = 1; platform_sprite[1][51][7] = 1; platform_sprite[1][51][8] = 1; platform_sprite[1][51][9] = 1; platform_sprite[1][51][20] = 1; platform_sprite[1][51][21] = 1; platform_sprite[1][51][22] = 1; platform_sprite[1][51][23] = 1; platform_sprite[1][51][24] = 1; platform_sprite[1][52][5] = 1; platform_sprite[1][52][6] = 1; platform_sprite[1][52][7] = 1; platform_sprite[1][52][8] = 1; platform_sprite[1][52][9] = 1; platform_sprite[1][52][20] = 1; platform_sprite[1][52][21] = 1; platform_sprite[1][52][22] = 1; platform_sprite[1][52][23] = 1; platform_sprite[1][52][24] = 1; platform_sprite[1][53][5] = 1; platform_sprite[1][53][6] = 1; platform_sprite[1][53][7] = 1; platform_sprite[1][53][8] = 1; platform_sprite[1][53][9] = 1; platform_sprite[1][53][20] = 1; platform_sprite[1][53][21] = 1; platform_sprite[1][53][22] = 1; platform_sprite[1][53][23] = 1; platform_sprite[1][53][24] = 1; platform_sprite[1][54][5] = 1; platform_sprite[1][54][6] = 1; platform_sprite[1][54][7] = 1; platform_sprite[1][54][8] = 1; platform_sprite[1][54][9] = 1; platform_sprite[1][54][20] = 1; platform_sprite[1][54][21] = 1; platform_sprite[1][54][22] = 1; platform_sprite[1][54][23] = 1; platform_sprite[1][54][24] = 1; platform_sprite[1][55][5] = 1; platform_sprite[1][55][6] = 1; platform_sprite[1][55][7] = 1; platform_sprite[1][55][8] = 1; platform_sprite[1][55][9] = 1; platform_sprite[1][55][20] = 1; platform_sprite[1][55][21] = 1; platform_sprite[1][55][22] = 1; platform_sprite[1][55][23] = 1; platform_sprite[1][55][24] = 1; platform_sprite[1][56][5] = 1; platform_sprite[1][56][6] = 1; platform_sprite[1][56][7] = 1; platform_sprite[1][56][8] = 1; platform_sprite[1][56][9] = 1; platform_sprite[1][56][20] = 1; platform_sprite[1][56][21] = 1; platform_sprite[1][56][22] = 1; platform_sprite[1][56][23] = 1; platform_sprite[1][56][24] = 1; platform_sprite[1][57][5] = 1; platform_sprite[1][57][6] = 1; platform_sprite[1][57][7] = 1; platform_sprite[1][57][8] = 1; platform_sprite[1][57][9] = 1; platform_sprite[1][57][20] = 1; platform_sprite[1][57][21] = 1; platform_sprite[1][57][22] = 1; platform_sprite[1][57][23] = 1; platform_sprite[1][57][24] = 1; platform_sprite[1][58][5] = 1; platform_sprite[1][58][6] = 1; platform_sprite[1][58][7] = 1; platform_sprite[1][58][8] = 1; platform_sprite[1][58][9] = 1; platform_sprite[1][58][20] = 1; platform_sprite[1][58][21] = 1; platform_sprite[1][58][22] = 1; platform_sprite[1][58][23] = 1; platform_sprite[1][58][24] = 1; platform_sprite[1][59][5] = 1; platform_sprite[1][59][6] = 1; platform_sprite[1][59][7] = 1; platform_sprite[1][59][8] = 1; platform_sprite[1][59][9] = 1; platform_sprite[1][59][20] = 1; platform_sprite[1][59][21] = 1; platform_sprite[1][59][22] = 1; platform_sprite[1][59][23] = 1; platform_sprite[1][59][24] = 1; platform_sprite[1][60][5] = 1; platform_sprite[1][60][6] = 1; platform_sprite[1][60][7] = 1; platform_sprite[1][60][8] = 1; platform_sprite[1][60][9] = 1; platform_sprite[1][60][20] = 1; platform_sprite[1][60][21] = 1; platform_sprite[1][60][22] = 1; platform_sprite[1][60][23] = 1; platform_sprite[1][60][24] = 1; platform_sprite[1][61][5] = 1; platform_sprite[1][61][6] = 1; platform_sprite[1][61][7] = 1; platform_sprite[1][61][8] = 1; platform_sprite[1][61][9] = 1; platform_sprite[1][61][20] = 1; platform_sprite[1][61][21] = 1; platform_sprite[1][61][22] = 1; platform_sprite[1][61][23] = 1; platform_sprite[1][61][24] = 1; platform_sprite[1][62][5] = 1; platform_sprite[1][62][6] = 1; platform_sprite[1][62][7] = 1; platform_sprite[1][62][8] = 1; platform_sprite[1][62][9] = 1; platform_sprite[1][62][20] = 1; platform_sprite[1][62][21] = 1; platform_sprite[1][62][22] = 1; platform_sprite[1][62][23] = 1; platform_sprite[1][62][24] = 1; platform_sprite[1][63][5] = 1; platform_sprite[1][63][6] = 1; platform_sprite[1][63][7] = 1; platform_sprite[1][63][8] = 1; platform_sprite[1][63][9] = 1; platform_sprite[1][63][20] = 1; platform_sprite[1][63][21] = 1; platform_sprite[1][63][22] = 1; platform_sprite[1][63][23] = 1; platform_sprite[1][63][24] = 1; platform_sprite[1][64][5] = 1; platform_sprite[1][64][6] = 1; platform_sprite[1][64][7] = 1; platform_sprite[1][64][8] = 1; platform_sprite[1][64][9] = 1; platform_sprite[1][64][20] = 1; platform_sprite[1][64][21] = 1; platform_sprite[1][64][22] = 1; platform_sprite[1][64][23] = 1; platform_sprite[1][64][24] = 1; platform_sprite[1][65][5] = 1; platform_sprite[1][65][6] = 1; platform_sprite[1][65][7] = 1; platform_sprite[1][65][8] = 1; platform_sprite[1][65][9] = 1; platform_sprite[1][65][20] = 1; platform_sprite[1][65][21] = 1; platform_sprite[1][65][22] = 1; platform_sprite[1][65][23] = 1; platform_sprite[1][65][24] = 1; platform_sprite[1][66][5] = 1; platform_sprite[1][66][6] = 1; platform_sprite[1][66][7] = 1; platform_sprite[1][66][8] = 1; platform_sprite[1][66][9] = 1; platform_sprite[1][66][20] = 1; platform_sprite[1][66][21] = 1; platform_sprite[1][66][22] = 1; platform_sprite[1][66][23] = 1; platform_sprite[1][66][24] = 1; platform_sprite[1][67][5] = 1; platform_sprite[1][67][6] = 1; platform_sprite[1][67][7] = 1; platform_sprite[1][67][8] = 1; platform_sprite[1][67][9] = 1; platform_sprite[1][67][20] = 1; platform_sprite[1][67][21] = 1; platform_sprite[1][67][22] = 1; platform_sprite[1][67][23] = 1; platform_sprite[1][67][24] = 1; platform_sprite[1][68][5] = 1; platform_sprite[1][68][6] = 1; platform_sprite[1][68][7] = 1; platform_sprite[1][68][8] = 1; platform_sprite[1][68][9] = 1; platform_sprite[1][68][20] = 1; platform_sprite[1][68][21] = 1; platform_sprite[1][68][22] = 1; platform_sprite[1][68][23] = 1; platform_sprite[1][68][24] = 1; platform_sprite[1][69][5] = 1; platform_sprite[1][69][6] = 1; platform_sprite[1][69][7] = 1; platform_sprite[1][69][8] = 1; platform_sprite[1][69][9] = 1; platform_sprite[1][69][20] = 1; platform_sprite[1][69][21] = 1; platform_sprite[1][69][22] = 1; platform_sprite[1][69][23] = 1; platform_sprite[1][69][24] = 1; platform_sprite[1][70][5] = 1; platform_sprite[1][70][6] = 1; platform_sprite[1][70][7] = 1; platform_sprite[1][70][8] = 1; platform_sprite[1][70][9] = 1; platform_sprite[1][70][20] = 1; platform_sprite[1][70][21] = 1; platform_sprite[1][70][22] = 1; platform_sprite[1][70][23] = 1; platform_sprite[1][70][24] = 1; platform_sprite[1][71][5] = 1; platform_sprite[1][71][6] = 1; platform_sprite[1][71][7] = 1; platform_sprite[1][71][8] = 1; platform_sprite[1][71][9] = 1; platform_sprite[1][71][20] = 1; platform_sprite[1][71][21] = 1; platform_sprite[1][71][22] = 1; platform_sprite[1][71][23] = 1; platform_sprite[1][71][24] = 1; platform_sprite[1][72][5] = 1; platform_sprite[1][72][6] = 1; platform_sprite[1][72][7] = 1; platform_sprite[1][72][8] = 1; platform_sprite[1][72][9] = 1; platform_sprite[1][72][20] = 1; platform_sprite[1][72][21] = 1; platform_sprite[1][72][22] = 1; platform_sprite[1][72][23] = 1; platform_sprite[1][72][24] = 1; platform_sprite[1][73][5] = 1; platform_sprite[1][73][6] = 1; platform_sprite[1][73][7] = 1; platform_sprite[1][73][8] = 1; platform_sprite[1][73][9] = 1; platform_sprite[1][73][20] = 1; platform_sprite[1][73][21] = 1; platform_sprite[1][73][22] = 1; platform_sprite[1][73][23] = 1; platform_sprite[1][73][24] = 1; platform_sprite[1][74][5] = 1; platform_sprite[1][74][6] = 1; platform_sprite[1][74][7] = 1; platform_sprite[1][74][8] = 1; platform_sprite[1][74][9] = 1; platform_sprite[1][74][20] = 1; platform_sprite[1][74][21] = 1; platform_sprite[1][74][22] = 1; platform_sprite[1][74][23] = 1; platform_sprite[1][74][24] = 1; platform_sprite[1][75][5] = 1; platform_sprite[1][75][6] = 1; platform_sprite[1][75][7] = 1; platform_sprite[1][75][8] = 1; platform_sprite[1][75][9] = 1; platform_sprite[1][75][20] = 1; platform_sprite[1][75][21] = 1; platform_sprite[1][75][22] = 1; platform_sprite[1][75][23] = 1; platform_sprite[1][75][24] = 1; platform_sprite[1][76][5] = 1; platform_sprite[1][76][6] = 1; platform_sprite[1][76][7] = 1; platform_sprite[1][76][8] = 1; platform_sprite[1][76][9] = 1; platform_sprite[1][76][20] = 1; platform_sprite[1][76][21] = 1; platform_sprite[1][76][22] = 1; platform_sprite[1][76][23] = 1; platform_sprite[1][76][24] = 1; platform_sprite[1][77][5] = 1; platform_sprite[1][77][6] = 1; platform_sprite[1][77][7] = 1; platform_sprite[1][77][8] = 1; platform_sprite[1][77][9] = 1; platform_sprite[1][77][20] = 1; platform_sprite[1][77][21] = 1; platform_sprite[1][77][22] = 1; platform_sprite[1][77][23] = 1; platform_sprite[1][77][24] = 1; platform_sprite[1][78][5] = 1; platform_sprite[1][78][6] = 1; platform_sprite[1][78][7] = 1; platform_sprite[1][78][8] = 1; platform_sprite[1][78][9] = 1; platform_sprite[1][78][20] = 1; platform_sprite[1][78][21] = 1; platform_sprite[1][78][22] = 1; platform_sprite[1][78][23] = 1; platform_sprite[1][78][24] = 1; platform_sprite[1][79][5] = 1; platform_sprite[1][79][6] = 1; platform_sprite[1][79][7] = 1; platform_sprite[1][79][8] = 1; platform_sprite[1][79][9] = 1; platform_sprite[1][79][20] = 1; platform_sprite[1][79][21] = 1; platform_sprite[1][79][22] = 1; platform_sprite[1][79][23] = 1; platform_sprite[1][79][24] = 1; platform_sprite[1][80][5] = 1; platform_sprite[1][80][6] = 1; platform_sprite[1][80][7] = 1; platform_sprite[1][80][8] = 1; platform_sprite[1][80][9] = 1; platform_sprite[1][80][20] = 1; platform_sprite[1][80][21] = 1; platform_sprite[1][80][22] = 1; platform_sprite[1][80][23] = 1; platform_sprite[1][80][24] = 1; platform_sprite[1][81][5] = 1; platform_sprite[1][81][6] = 1; platform_sprite[1][81][7] = 1; platform_sprite[1][81][8] = 1; platform_sprite[1][81][9] = 1; platform_sprite[1][81][20] = 1; platform_sprite[1][81][21] = 1; platform_sprite[1][81][22] = 1; platform_sprite[1][81][23] = 1; platform_sprite[1][81][24] = 1; platform_sprite[1][82][5] = 1; platform_sprite[1][82][6] = 1; platform_sprite[1][82][7] = 1; platform_sprite[1][82][8] = 1; platform_sprite[1][82][9] = 1; platform_sprite[1][82][20] = 1; platform_sprite[1][82][21] = 1; platform_sprite[1][82][22] = 1; platform_sprite[1][82][23] = 1; platform_sprite[1][82][24] = 1; platform_sprite[1][83][5] = 1; platform_sprite[1][83][6] = 1; platform_sprite[1][83][7] = 1; platform_sprite[1][83][8] = 1; platform_sprite[1][83][9] = 1; platform_sprite[1][83][20] = 1; platform_sprite[1][83][21] = 1; platform_sprite[1][83][22] = 1; platform_sprite[1][83][23] = 1; platform_sprite[1][83][24] = 1; platform_sprite[1][84][5] = 1; platform_sprite[1][84][6] = 1; platform_sprite[1][84][7] = 1; platform_sprite[1][84][8] = 1; platform_sprite[1][84][9] = 1; platform_sprite[1][84][20] = 1; platform_sprite[1][84][21] = 1; platform_sprite[1][84][22] = 1; platform_sprite[1][84][23] = 1; platform_sprite[1][84][24] = 1; platform_sprite[1][85][5] = 1; platform_sprite[1][85][6] = 1; platform_sprite[1][85][7] = 1; platform_sprite[1][85][8] = 1; platform_sprite[1][85][9] = 1; platform_sprite[1][85][20] = 1; platform_sprite[1][85][21] = 1; platform_sprite[1][85][22] = 1; platform_sprite[1][85][23] = 1; platform_sprite[1][85][24] = 1; platform_sprite[1][86][5] = 1; platform_sprite[1][86][6] = 1; platform_sprite[1][86][7] = 1; platform_sprite[1][86][8] = 1; platform_sprite[1][86][9] = 1; platform_sprite[1][86][20] = 1; platform_sprite[1][86][21] = 1; platform_sprite[1][86][22] = 1; platform_sprite[1][86][23] = 1; platform_sprite[1][86][24] = 1; platform_sprite[1][87][5] = 1; platform_sprite[1][87][6] = 1; platform_sprite[1][87][7] = 1; platform_sprite[1][87][8] = 1; platform_sprite[1][87][9] = 1; platform_sprite[1][87][20] = 1; platform_sprite[1][87][21] = 1; platform_sprite[1][87][22] = 1; platform_sprite[1][87][23] = 1; platform_sprite[1][87][24] = 1; platform_sprite[1][88][5] = 1; platform_sprite[1][88][6] = 1; platform_sprite[1][88][7] = 1; platform_sprite[1][88][8] = 1; platform_sprite[1][88][9] = 1; platform_sprite[1][88][20] = 1; platform_sprite[1][88][21] = 1; platform_sprite[1][88][22] = 1; platform_sprite[1][88][23] = 1; platform_sprite[1][88][24] = 1; platform_sprite[1][89][5] = 1; platform_sprite[1][89][6] = 1; platform_sprite[1][89][7] = 1; platform_sprite[1][89][8] = 1; platform_sprite[1][89][9] = 1; platform_sprite[1][89][20] = 1; platform_sprite[1][89][21] = 1; platform_sprite[1][89][22] = 1; platform_sprite[1][89][23] = 1; platform_sprite[1][89][24] = 1; platform_sprite[1][90][10] = 1; platform_sprite[1][90][11] = 1; platform_sprite[1][90][12] = 1; platform_sprite[1][90][13] = 1; platform_sprite[1][90][14] = 1; platform_sprite[1][90][15] = 1; platform_sprite[1][90][16] = 1; platform_sprite[1][90][17] = 1; platform_sprite[1][90][18] = 1; platform_sprite[1][90][19] = 1; platform_sprite[1][91][10] = 1; platform_sprite[1][91][11] = 1; platform_sprite[1][91][12] = 1; platform_sprite[1][91][13] = 1; platform_sprite[1][91][14] = 1; platform_sprite[1][91][15] = 1; platform_sprite[1][91][16] = 1; platform_sprite[1][91][17] = 1; platform_sprite[1][91][18] = 1; platform_sprite[1][91][19] = 1; platform_sprite[1][92][10] = 1; platform_sprite[1][92][11] = 1; platform_sprite[1][92][12] = 1; platform_sprite[1][92][13] = 1; platform_sprite[1][92][14] = 1; platform_sprite[1][92][15] = 1; platform_sprite[1][92][16] = 1; platform_sprite[1][92][17] = 1; platform_sprite[1][92][18] = 1; platform_sprite[1][92][19] = 1; platform_sprite[1][93][10] = 1; platform_sprite[1][93][11] = 1; platform_sprite[1][93][12] = 1; platform_sprite[1][93][13] = 1; platform_sprite[1][93][14] = 1; platform_sprite[1][93][15] = 1; platform_sprite[1][93][16] = 1; platform_sprite[1][93][17] = 1; platform_sprite[1][93][18] = 1; platform_sprite[1][93][19] = 1; platform_sprite[1][94][10] = 1; platform_sprite[1][94][11] = 1; platform_sprite[1][94][12] = 1; platform_sprite[1][94][13] = 1; platform_sprite[1][94][14] = 1; platform_sprite[1][94][15] = 1; platform_sprite[1][94][16] = 1; platform_sprite[1][94][17] = 1; platform_sprite[1][94][18] = 1; platform_sprite[1][94][19] = 1; 
					platform_sprite[2][5][10] = 1; platform_sprite[2][5][11] = 1; platform_sprite[2][5][12] = 1; platform_sprite[2][5][13] = 1; platform_sprite[2][5][14] = 1; platform_sprite[2][5][15] = 1; platform_sprite[2][5][16] = 1; platform_sprite[2][5][17] = 1; platform_sprite[2][5][18] = 1; platform_sprite[2][5][19] = 1; platform_sprite[2][6][10] = 1; platform_sprite[2][6][11] = 1; platform_sprite[2][6][12] = 1; platform_sprite[2][6][13] = 1; platform_sprite[2][6][14] = 1; platform_sprite[2][6][15] = 1; platform_sprite[2][6][16] = 1; platform_sprite[2][6][17] = 1; platform_sprite[2][6][18] = 1; platform_sprite[2][6][19] = 1; platform_sprite[2][7][10] = 1; platform_sprite[2][7][11] = 1; platform_sprite[2][7][12] = 1; platform_sprite[2][7][13] = 1; platform_sprite[2][7][14] = 1; platform_sprite[2][7][15] = 1; platform_sprite[2][7][16] = 1; platform_sprite[2][7][17] = 1; platform_sprite[2][7][18] = 1; platform_sprite[2][7][19] = 1; platform_sprite[2][8][10] = 1; platform_sprite[2][8][11] = 1; platform_sprite[2][8][12] = 1; platform_sprite[2][8][13] = 1; platform_sprite[2][8][14] = 1; platform_sprite[2][8][15] = 1; platform_sprite[2][8][16] = 1; platform_sprite[2][8][17] = 1; platform_sprite[2][8][18] = 1; platform_sprite[2][8][19] = 1; platform_sprite[2][9][10] = 1; platform_sprite[2][9][11] = 1; platform_sprite[2][9][12] = 1; platform_sprite[2][9][13] = 1; platform_sprite[2][9][14] = 1; platform_sprite[2][9][15] = 1; platform_sprite[2][9][16] = 1; platform_sprite[2][9][17] = 1; platform_sprite[2][9][18] = 1; platform_sprite[2][9][19] = 1; platform_sprite[2][9][20] = 1; platform_sprite[2][9][21] = 1; platform_sprite[2][9][22] = 1; platform_sprite[2][9][23] = 1; platform_sprite[2][9][24] = 1; platform_sprite[2][10][5] = 1; platform_sprite[2][10][6] = 1; platform_sprite[2][10][7] = 1; platform_sprite[2][10][8] = 1; platform_sprite[2][10][9] = 1; platform_sprite[2][10][20] = 1; platform_sprite[2][10][21] = 1; platform_sprite[2][10][22] = 1; platform_sprite[2][10][23] = 1; platform_sprite[2][10][24] = 1; platform_sprite[2][11][5] = 1; platform_sprite[2][11][6] = 1; platform_sprite[2][11][7] = 1; platform_sprite[2][11][8] = 1; platform_sprite[2][11][9] = 1; platform_sprite[2][11][20] = 1; platform_sprite[2][11][21] = 1; platform_sprite[2][11][22] = 1; platform_sprite[2][11][23] = 1; platform_sprite[2][11][24] = 1; platform_sprite[2][12][5] = 1; platform_sprite[2][12][6] = 1; platform_sprite[2][12][7] = 1; platform_sprite[2][12][8] = 1; platform_sprite[2][12][9] = 1; platform_sprite[2][12][20] = 1; platform_sprite[2][12][21] = 1; platform_sprite[2][12][22] = 1; platform_sprite[2][12][23] = 1; platform_sprite[2][12][24] = 1; platform_sprite[2][13][5] = 1; platform_sprite[2][13][6] = 1; platform_sprite[2][13][7] = 1; platform_sprite[2][13][8] = 1; platform_sprite[2][13][9] = 1; platform_sprite[2][13][20] = 1; platform_sprite[2][13][21] = 1; platform_sprite[2][13][22] = 1; platform_sprite[2][13][23] = 1; platform_sprite[2][13][24] = 1; platform_sprite[2][14][5] = 1; platform_sprite[2][14][6] = 1; platform_sprite[2][14][7] = 1; platform_sprite[2][14][8] = 1; platform_sprite[2][14][9] = 1; platform_sprite[2][14][20] = 1; platform_sprite[2][14][21] = 1; platform_sprite[2][14][22] = 1; platform_sprite[2][14][23] = 1; platform_sprite[2][14][24] = 1; platform_sprite[2][15][5] = 1; platform_sprite[2][15][6] = 1; platform_sprite[2][15][7] = 1; platform_sprite[2][15][8] = 1; platform_sprite[2][15][9] = 1; platform_sprite[2][15][20] = 1; platform_sprite[2][15][21] = 1; platform_sprite[2][15][22] = 1; platform_sprite[2][15][23] = 1; platform_sprite[2][15][24] = 1; platform_sprite[2][16][5] = 1; platform_sprite[2][16][6] = 1; platform_sprite[2][16][7] = 1; platform_sprite[2][16][8] = 1; platform_sprite[2][16][9] = 1; platform_sprite[2][16][20] = 1; platform_sprite[2][16][21] = 1; platform_sprite[2][16][22] = 1; platform_sprite[2][16][23] = 1; platform_sprite[2][16][24] = 1; platform_sprite[2][17][5] = 1; platform_sprite[2][17][6] = 1; platform_sprite[2][17][7] = 1; platform_sprite[2][17][8] = 1; platform_sprite[2][17][9] = 1; platform_sprite[2][17][20] = 1; platform_sprite[2][17][21] = 1; platform_sprite[2][17][22] = 1; platform_sprite[2][17][23] = 1; platform_sprite[2][17][24] = 1; platform_sprite[2][18][5] = 1; platform_sprite[2][18][6] = 1; platform_sprite[2][18][7] = 1; platform_sprite[2][18][8] = 1; platform_sprite[2][18][9] = 1; platform_sprite[2][18][20] = 1; platform_sprite[2][18][21] = 1; platform_sprite[2][18][22] = 1; platform_sprite[2][18][23] = 1; platform_sprite[2][18][24] = 1; platform_sprite[2][19][5] = 1; platform_sprite[2][19][6] = 1; platform_sprite[2][19][7] = 1; platform_sprite[2][19][8] = 1; platform_sprite[2][19][9] = 1; platform_sprite[2][19][20] = 1; platform_sprite[2][19][21] = 1; platform_sprite[2][19][22] = 1; platform_sprite[2][19][23] = 1; platform_sprite[2][19][24] = 1; platform_sprite[2][20][5] = 1; platform_sprite[2][20][6] = 1; platform_sprite[2][20][7] = 1; platform_sprite[2][20][8] = 1; platform_sprite[2][20][9] = 1; platform_sprite[2][20][20] = 1; platform_sprite[2][20][21] = 1; platform_sprite[2][20][22] = 1; platform_sprite[2][20][23] = 1; platform_sprite[2][20][24] = 1; platform_sprite[2][21][5] = 1; platform_sprite[2][21][6] = 1; platform_sprite[2][21][7] = 1; platform_sprite[2][21][8] = 1; platform_sprite[2][21][9] = 1; platform_sprite[2][21][20] = 1; platform_sprite[2][21][21] = 1; platform_sprite[2][21][22] = 1; platform_sprite[2][21][23] = 1; platform_sprite[2][21][24] = 1; platform_sprite[2][22][5] = 1; platform_sprite[2][22][6] = 1; platform_sprite[2][22][7] = 1; platform_sprite[2][22][8] = 1; platform_sprite[2][22][9] = 1; platform_sprite[2][22][20] = 1; platform_sprite[2][22][21] = 1; platform_sprite[2][22][22] = 1; platform_sprite[2][22][23] = 1; platform_sprite[2][22][24] = 1; platform_sprite[2][23][5] = 1; platform_sprite[2][23][6] = 1; platform_sprite[2][23][7] = 1; platform_sprite[2][23][8] = 1; platform_sprite[2][23][9] = 1; platform_sprite[2][23][20] = 1; platform_sprite[2][23][21] = 1; platform_sprite[2][23][22] = 1; platform_sprite[2][23][23] = 1; platform_sprite[2][23][24] = 1; platform_sprite[2][24][5] = 1; platform_sprite[2][24][6] = 1; platform_sprite[2][24][7] = 1; platform_sprite[2][24][8] = 1; platform_sprite[2][24][9] = 1; platform_sprite[2][24][20] = 1; platform_sprite[2][24][21] = 1; platform_sprite[2][24][22] = 1; platform_sprite[2][24][23] = 1; platform_sprite[2][24][24] = 1; platform_sprite[2][25][5] = 1; platform_sprite[2][25][6] = 1; platform_sprite[2][25][7] = 1; platform_sprite[2][25][8] = 1; platform_sprite[2][25][9] = 1; platform_sprite[2][25][20] = 1; platform_sprite[2][25][21] = 1; platform_sprite[2][25][22] = 1; platform_sprite[2][25][23] = 1; platform_sprite[2][25][24] = 1; platform_sprite[2][26][5] = 1; platform_sprite[2][26][6] = 1; platform_sprite[2][26][7] = 1; platform_sprite[2][26][8] = 1; platform_sprite[2][26][9] = 1; platform_sprite[2][26][20] = 1; platform_sprite[2][26][21] = 1; platform_sprite[2][26][22] = 1; platform_sprite[2][26][23] = 1; platform_sprite[2][26][24] = 1; platform_sprite[2][27][5] = 1; platform_sprite[2][27][6] = 1; platform_sprite[2][27][7] = 1; platform_sprite[2][27][8] = 1; platform_sprite[2][27][9] = 1; platform_sprite[2][27][20] = 1; platform_sprite[2][27][21] = 1; platform_sprite[2][27][22] = 1; platform_sprite[2][27][23] = 1; platform_sprite[2][27][24] = 1; platform_sprite[2][28][5] = 1; platform_sprite[2][28][6] = 1; platform_sprite[2][28][7] = 1; platform_sprite[2][28][8] = 1; platform_sprite[2][28][9] = 1; platform_sprite[2][28][20] = 1; platform_sprite[2][28][21] = 1; platform_sprite[2][28][22] = 1; platform_sprite[2][28][23] = 1; platform_sprite[2][28][24] = 1; platform_sprite[2][29][5] = 1; platform_sprite[2][29][6] = 1; platform_sprite[2][29][7] = 1; platform_sprite[2][29][8] = 1; platform_sprite[2][29][9] = 1; platform_sprite[2][29][20] = 1; platform_sprite[2][29][21] = 1; platform_sprite[2][29][22] = 1; platform_sprite[2][29][23] = 1; platform_sprite[2][29][24] = 1; platform_sprite[2][30][5] = 1; platform_sprite[2][30][6] = 1; platform_sprite[2][30][7] = 1; platform_sprite[2][30][8] = 1; platform_sprite[2][30][9] = 1; platform_sprite[2][30][20] = 1; platform_sprite[2][30][21] = 1; platform_sprite[2][30][22] = 1; platform_sprite[2][30][23] = 1; platform_sprite[2][30][24] = 1; platform_sprite[2][31][5] = 1; platform_sprite[2][31][6] = 1; platform_sprite[2][31][7] = 1; platform_sprite[2][31][8] = 1; platform_sprite[2][31][9] = 1; platform_sprite[2][31][20] = 1; platform_sprite[2][31][21] = 1; platform_sprite[2][31][22] = 1; platform_sprite[2][31][23] = 1; platform_sprite[2][31][24] = 1; platform_sprite[2][32][5] = 1; platform_sprite[2][32][6] = 1; platform_sprite[2][32][7] = 1; platform_sprite[2][32][8] = 1; platform_sprite[2][32][9] = 1; platform_sprite[2][32][20] = 1; platform_sprite[2][32][21] = 1; platform_sprite[2][32][22] = 1; platform_sprite[2][32][23] = 1; platform_sprite[2][32][24] = 1; platform_sprite[2][33][5] = 1; platform_sprite[2][33][6] = 1; platform_sprite[2][33][7] = 1; platform_sprite[2][33][8] = 1; platform_sprite[2][33][9] = 1; platform_sprite[2][33][20] = 1; platform_sprite[2][33][21] = 1; platform_sprite[2][33][22] = 1; platform_sprite[2][33][23] = 1; platform_sprite[2][33][24] = 1; platform_sprite[2][34][5] = 1; platform_sprite[2][34][6] = 1; platform_sprite[2][34][7] = 1; platform_sprite[2][34][8] = 1; platform_sprite[2][34][9] = 1; platform_sprite[2][34][20] = 1; platform_sprite[2][34][21] = 1; platform_sprite[2][34][22] = 1; platform_sprite[2][34][23] = 1; platform_sprite[2][34][24] = 1; platform_sprite[2][35][5] = 1; platform_sprite[2][35][6] = 1; platform_sprite[2][35][7] = 1; platform_sprite[2][35][8] = 1; platform_sprite[2][35][9] = 1; platform_sprite[2][35][20] = 1; platform_sprite[2][35][21] = 1; platform_sprite[2][35][22] = 1; platform_sprite[2][35][23] = 1; platform_sprite[2][35][24] = 1; platform_sprite[2][36][5] = 1; platform_sprite[2][36][6] = 1; platform_sprite[2][36][7] = 1; platform_sprite[2][36][8] = 1; platform_sprite[2][36][9] = 1; platform_sprite[2][36][20] = 1; platform_sprite[2][36][21] = 1; platform_sprite[2][36][22] = 1; platform_sprite[2][36][23] = 1; platform_sprite[2][36][24] = 1; platform_sprite[2][37][5] = 1; platform_sprite[2][37][6] = 1; platform_sprite[2][37][7] = 1; platform_sprite[2][37][8] = 1; platform_sprite[2][37][9] = 1; platform_sprite[2][37][20] = 1; platform_sprite[2][37][21] = 1; platform_sprite[2][37][22] = 1; platform_sprite[2][37][23] = 1; platform_sprite[2][37][24] = 1; platform_sprite[2][38][5] = 1; platform_sprite[2][38][6] = 1; platform_sprite[2][38][7] = 1; platform_sprite[2][38][8] = 1; platform_sprite[2][38][9] = 1; platform_sprite[2][38][20] = 1; platform_sprite[2][38][21] = 1; platform_sprite[2][38][22] = 1; platform_sprite[2][38][23] = 1; platform_sprite[2][38][24] = 1; platform_sprite[2][39][5] = 1; platform_sprite[2][39][6] = 1; platform_sprite[2][39][7] = 1; platform_sprite[2][39][8] = 1; platform_sprite[2][39][9] = 1; platform_sprite[2][39][20] = 1; platform_sprite[2][39][21] = 1; platform_sprite[2][39][22] = 1; platform_sprite[2][39][23] = 1; platform_sprite[2][39][24] = 1; platform_sprite[2][40][5] = 1; platform_sprite[2][40][6] = 1; platform_sprite[2][40][7] = 1; platform_sprite[2][40][8] = 1; platform_sprite[2][40][9] = 1; platform_sprite[2][40][20] = 1; platform_sprite[2][40][21] = 1; platform_sprite[2][40][22] = 1; platform_sprite[2][40][23] = 1; platform_sprite[2][40][24] = 1; platform_sprite[2][41][5] = 1; platform_sprite[2][41][6] = 1; platform_sprite[2][41][7] = 1; platform_sprite[2][41][8] = 1; platform_sprite[2][41][9] = 1; platform_sprite[2][41][20] = 1; platform_sprite[2][41][21] = 1; platform_sprite[2][41][22] = 1; platform_sprite[2][41][23] = 1; platform_sprite[2][41][24] = 1; platform_sprite[2][42][5] = 1; platform_sprite[2][42][6] = 1; platform_sprite[2][42][7] = 1; platform_sprite[2][42][8] = 1; platform_sprite[2][42][9] = 1; platform_sprite[2][42][20] = 1; platform_sprite[2][42][21] = 1; platform_sprite[2][42][22] = 1; platform_sprite[2][42][23] = 1; platform_sprite[2][42][24] = 1; platform_sprite[2][43][5] = 1; platform_sprite[2][43][6] = 1; platform_sprite[2][43][7] = 1; platform_sprite[2][43][8] = 1; platform_sprite[2][43][9] = 1; platform_sprite[2][43][20] = 1; platform_sprite[2][43][21] = 1; platform_sprite[2][43][22] = 1; platform_sprite[2][43][23] = 1; platform_sprite[2][43][24] = 1; platform_sprite[2][44][5] = 1; platform_sprite[2][44][6] = 1; platform_sprite[2][44][7] = 1; platform_sprite[2][44][8] = 1; platform_sprite[2][44][9] = 1; platform_sprite[2][44][20] = 1; platform_sprite[2][44][21] = 1; platform_sprite[2][44][22] = 1; platform_sprite[2][44][23] = 1; platform_sprite[2][44][24] = 1; platform_sprite[2][45][5] = 1; platform_sprite[2][45][6] = 1; platform_sprite[2][45][7] = 1; platform_sprite[2][45][8] = 1; platform_sprite[2][45][9] = 1; platform_sprite[2][45][20] = 1; platform_sprite[2][45][21] = 1; platform_sprite[2][45][22] = 1; platform_sprite[2][45][23] = 1; platform_sprite[2][45][24] = 1; platform_sprite[2][46][5] = 1; platform_sprite[2][46][6] = 1; platform_sprite[2][46][7] = 1; platform_sprite[2][46][8] = 1; platform_sprite[2][46][9] = 1; platform_sprite[2][46][20] = 1; platform_sprite[2][46][21] = 1; platform_sprite[2][46][22] = 1; platform_sprite[2][46][23] = 1; platform_sprite[2][46][24] = 1; platform_sprite[2][47][5] = 1; platform_sprite[2][47][6] = 1; platform_sprite[2][47][7] = 1; platform_sprite[2][47][8] = 1; platform_sprite[2][47][9] = 1; platform_sprite[2][47][20] = 1; platform_sprite[2][47][21] = 1; platform_sprite[2][47][22] = 1; platform_sprite[2][47][23] = 1; platform_sprite[2][47][24] = 1; platform_sprite[2][48][5] = 1; platform_sprite[2][48][6] = 1; platform_sprite[2][48][7] = 1; platform_sprite[2][48][8] = 1; platform_sprite[2][48][9] = 1; platform_sprite[2][48][20] = 1; platform_sprite[2][48][21] = 1; platform_sprite[2][48][22] = 1; platform_sprite[2][48][23] = 1; platform_sprite[2][48][24] = 1; platform_sprite[2][49][5] = 1; platform_sprite[2][49][6] = 1; platform_sprite[2][49][7] = 1; platform_sprite[2][49][8] = 1; platform_sprite[2][49][9] = 1; platform_sprite[2][49][20] = 1; platform_sprite[2][49][21] = 1; platform_sprite[2][49][22] = 1; platform_sprite[2][49][23] = 1; platform_sprite[2][49][24] = 1; platform_sprite[2][50][5] = 1; platform_sprite[2][50][6] = 1; platform_sprite[2][50][7] = 1; platform_sprite[2][50][8] = 1; platform_sprite[2][50][9] = 1; platform_sprite[2][50][20] = 1; platform_sprite[2][50][21] = 1; platform_sprite[2][50][22] = 1; platform_sprite[2][50][23] = 1; platform_sprite[2][50][24] = 1; platform_sprite[2][51][5] = 1; platform_sprite[2][51][6] = 1; platform_sprite[2][51][7] = 1; platform_sprite[2][51][8] = 1; platform_sprite[2][51][9] = 1; platform_sprite[2][51][20] = 1; platform_sprite[2][51][21] = 1; platform_sprite[2][51][22] = 1; platform_sprite[2][51][23] = 1; platform_sprite[2][51][24] = 1; platform_sprite[2][52][5] = 1; platform_sprite[2][52][6] = 1; platform_sprite[2][52][7] = 1; platform_sprite[2][52][8] = 1; platform_sprite[2][52][9] = 1; platform_sprite[2][52][20] = 1; platform_sprite[2][52][21] = 1; platform_sprite[2][52][22] = 1; platform_sprite[2][52][23] = 1; platform_sprite[2][52][24] = 1; platform_sprite[2][53][5] = 1; platform_sprite[2][53][6] = 1; platform_sprite[2][53][7] = 1; platform_sprite[2][53][8] = 1; platform_sprite[2][53][9] = 1; platform_sprite[2][53][20] = 1; platform_sprite[2][53][21] = 1; platform_sprite[2][53][22] = 1; platform_sprite[2][53][23] = 1; platform_sprite[2][53][24] = 1; platform_sprite[2][54][5] = 1; platform_sprite[2][54][6] = 1; platform_sprite[2][54][7] = 1; platform_sprite[2][54][8] = 1; platform_sprite[2][54][9] = 1; platform_sprite[2][54][20] = 1; platform_sprite[2][54][21] = 1; platform_sprite[2][54][22] = 1; platform_sprite[2][54][23] = 1; platform_sprite[2][54][24] = 1; platform_sprite[2][55][5] = 1; platform_sprite[2][55][6] = 1; platform_sprite[2][55][7] = 1; platform_sprite[2][55][8] = 1; platform_sprite[2][55][9] = 1; platform_sprite[2][55][20] = 1; platform_sprite[2][55][21] = 1; platform_sprite[2][55][22] = 1; platform_sprite[2][55][23] = 1; platform_sprite[2][55][24] = 1; platform_sprite[2][56][5] = 1; platform_sprite[2][56][6] = 1; platform_sprite[2][56][7] = 1; platform_sprite[2][56][8] = 1; platform_sprite[2][56][9] = 1; platform_sprite[2][56][20] = 1; platform_sprite[2][56][21] = 1; platform_sprite[2][56][22] = 1; platform_sprite[2][56][23] = 1; platform_sprite[2][56][24] = 1; platform_sprite[2][57][5] = 1; platform_sprite[2][57][6] = 1; platform_sprite[2][57][7] = 1; platform_sprite[2][57][8] = 1; platform_sprite[2][57][9] = 1; platform_sprite[2][57][20] = 1; platform_sprite[2][57][21] = 1; platform_sprite[2][57][22] = 1; platform_sprite[2][57][23] = 1; platform_sprite[2][57][24] = 1; platform_sprite[2][58][5] = 1; platform_sprite[2][58][6] = 1; platform_sprite[2][58][7] = 1; platform_sprite[2][58][8] = 1; platform_sprite[2][58][9] = 1; platform_sprite[2][58][20] = 1; platform_sprite[2][58][21] = 1; platform_sprite[2][58][22] = 1; platform_sprite[2][58][23] = 1; platform_sprite[2][58][24] = 1; platform_sprite[2][59][5] = 1; platform_sprite[2][59][6] = 1; platform_sprite[2][59][7] = 1; platform_sprite[2][59][8] = 1; platform_sprite[2][59][9] = 1; platform_sprite[2][59][20] = 1; platform_sprite[2][59][21] = 1; platform_sprite[2][59][22] = 1; platform_sprite[2][59][23] = 1; platform_sprite[2][59][24] = 1; platform_sprite[2][60][5] = 1; platform_sprite[2][60][6] = 1; platform_sprite[2][60][7] = 1; platform_sprite[2][60][8] = 1; platform_sprite[2][60][9] = 1; platform_sprite[2][60][20] = 1; platform_sprite[2][60][21] = 1; platform_sprite[2][60][22] = 1; platform_sprite[2][60][23] = 1; platform_sprite[2][60][24] = 1; platform_sprite[2][61][5] = 1; platform_sprite[2][61][6] = 1; platform_sprite[2][61][7] = 1; platform_sprite[2][61][8] = 1; platform_sprite[2][61][9] = 1; platform_sprite[2][61][20] = 1; platform_sprite[2][61][21] = 1; platform_sprite[2][61][22] = 1; platform_sprite[2][61][23] = 1; platform_sprite[2][61][24] = 1; platform_sprite[2][62][5] = 1; platform_sprite[2][62][6] = 1; platform_sprite[2][62][7] = 1; platform_sprite[2][62][8] = 1; platform_sprite[2][62][9] = 1; platform_sprite[2][62][20] = 1; platform_sprite[2][62][21] = 1; platform_sprite[2][62][22] = 1; platform_sprite[2][62][23] = 1; platform_sprite[2][62][24] = 1; platform_sprite[2][63][5] = 1; platform_sprite[2][63][6] = 1; platform_sprite[2][63][7] = 1; platform_sprite[2][63][8] = 1; platform_sprite[2][63][9] = 1; platform_sprite[2][63][20] = 1; platform_sprite[2][63][21] = 1; platform_sprite[2][63][22] = 1; platform_sprite[2][63][23] = 1; platform_sprite[2][63][24] = 1; platform_sprite[2][64][5] = 1; platform_sprite[2][64][6] = 1; platform_sprite[2][64][7] = 1; platform_sprite[2][64][8] = 1; platform_sprite[2][64][9] = 1; platform_sprite[2][64][20] = 1; platform_sprite[2][64][21] = 1; platform_sprite[2][64][22] = 1; platform_sprite[2][64][23] = 1; platform_sprite[2][64][24] = 1; platform_sprite[2][65][5] = 1; platform_sprite[2][65][6] = 1; platform_sprite[2][65][7] = 1; platform_sprite[2][65][8] = 1; platform_sprite[2][65][9] = 1; platform_sprite[2][65][20] = 1; platform_sprite[2][65][21] = 1; platform_sprite[2][65][22] = 1; platform_sprite[2][65][23] = 1; platform_sprite[2][65][24] = 1; platform_sprite[2][66][5] = 1; platform_sprite[2][66][6] = 1; platform_sprite[2][66][7] = 1; platform_sprite[2][66][8] = 1; platform_sprite[2][66][9] = 1; platform_sprite[2][66][20] = 1; platform_sprite[2][66][21] = 1; platform_sprite[2][66][22] = 1; platform_sprite[2][66][23] = 1; platform_sprite[2][66][24] = 1; platform_sprite[2][67][5] = 1; platform_sprite[2][67][6] = 1; platform_sprite[2][67][7] = 1; platform_sprite[2][67][8] = 1; platform_sprite[2][67][9] = 1; platform_sprite[2][67][20] = 1; platform_sprite[2][67][21] = 1; platform_sprite[2][67][22] = 1; platform_sprite[2][67][23] = 1; platform_sprite[2][67][24] = 1; platform_sprite[2][68][5] = 1; platform_sprite[2][68][6] = 1; platform_sprite[2][68][7] = 1; platform_sprite[2][68][8] = 1; platform_sprite[2][68][9] = 1; platform_sprite[2][68][20] = 1; platform_sprite[2][68][21] = 1; platform_sprite[2][68][22] = 1; platform_sprite[2][68][23] = 1; platform_sprite[2][68][24] = 1; platform_sprite[2][69][5] = 1; platform_sprite[2][69][6] = 1; platform_sprite[2][69][7] = 1; platform_sprite[2][69][8] = 1; platform_sprite[2][69][9] = 1; platform_sprite[2][69][20] = 1; platform_sprite[2][69][21] = 1; platform_sprite[2][69][22] = 1; platform_sprite[2][69][23] = 1; platform_sprite[2][69][24] = 1; platform_sprite[2][70][5] = 1; platform_sprite[2][70][6] = 1; platform_sprite[2][70][7] = 1; platform_sprite[2][70][8] = 1; platform_sprite[2][70][9] = 1; platform_sprite[2][70][20] = 1; platform_sprite[2][70][21] = 1; platform_sprite[2][70][22] = 1; platform_sprite[2][70][23] = 1; platform_sprite[2][70][24] = 1; platform_sprite[2][71][5] = 1; platform_sprite[2][71][6] = 1; platform_sprite[2][71][7] = 1; platform_sprite[2][71][8] = 1; platform_sprite[2][71][9] = 1; platform_sprite[2][71][20] = 1; platform_sprite[2][71][21] = 1; platform_sprite[2][71][22] = 1; platform_sprite[2][71][23] = 1; platform_sprite[2][71][24] = 1; platform_sprite[2][72][5] = 1; platform_sprite[2][72][6] = 1; platform_sprite[2][72][7] = 1; platform_sprite[2][72][8] = 1; platform_sprite[2][72][9] = 1; platform_sprite[2][72][20] = 1; platform_sprite[2][72][21] = 1; platform_sprite[2][72][22] = 1; platform_sprite[2][72][23] = 1; platform_sprite[2][72][24] = 1; platform_sprite[2][73][5] = 1; platform_sprite[2][73][6] = 1; platform_sprite[2][73][7] = 1; platform_sprite[2][73][8] = 1; platform_sprite[2][73][9] = 1; platform_sprite[2][73][20] = 1; platform_sprite[2][73][21] = 1; platform_sprite[2][73][22] = 1; platform_sprite[2][73][23] = 1; platform_sprite[2][73][24] = 1; platform_sprite[2][74][5] = 1; platform_sprite[2][74][6] = 1; platform_sprite[2][74][7] = 1; platform_sprite[2][74][8] = 1; platform_sprite[2][74][9] = 1; platform_sprite[2][74][20] = 1; platform_sprite[2][74][21] = 1; platform_sprite[2][74][22] = 1; platform_sprite[2][74][23] = 1; platform_sprite[2][74][24] = 1; platform_sprite[2][75][5] = 1; platform_sprite[2][75][6] = 1; platform_sprite[2][75][7] = 1; platform_sprite[2][75][8] = 1; platform_sprite[2][75][9] = 1; platform_sprite[2][75][20] = 1; platform_sprite[2][75][21] = 1; platform_sprite[2][75][22] = 1; platform_sprite[2][75][23] = 1; platform_sprite[2][75][24] = 1; platform_sprite[2][76][5] = 1; platform_sprite[2][76][6] = 1; platform_sprite[2][76][7] = 1; platform_sprite[2][76][8] = 1; platform_sprite[2][76][9] = 1; platform_sprite[2][76][20] = 1; platform_sprite[2][76][21] = 1; platform_sprite[2][76][22] = 1; platform_sprite[2][76][23] = 1; platform_sprite[2][76][24] = 1; platform_sprite[2][77][5] = 1; platform_sprite[2][77][6] = 1; platform_sprite[2][77][7] = 1; platform_sprite[2][77][8] = 1; platform_sprite[2][77][9] = 1; platform_sprite[2][77][20] = 1; platform_sprite[2][77][21] = 1; platform_sprite[2][77][22] = 1; platform_sprite[2][77][23] = 1; platform_sprite[2][77][24] = 1; platform_sprite[2][78][5] = 1; platform_sprite[2][78][6] = 1; platform_sprite[2][78][7] = 1; platform_sprite[2][78][8] = 1; platform_sprite[2][78][9] = 1; platform_sprite[2][78][20] = 1; platform_sprite[2][78][21] = 1; platform_sprite[2][78][22] = 1; platform_sprite[2][78][23] = 1; platform_sprite[2][78][24] = 1; platform_sprite[2][79][5] = 1; platform_sprite[2][79][6] = 1; platform_sprite[2][79][7] = 1; platform_sprite[2][79][8] = 1; platform_sprite[2][79][9] = 1; platform_sprite[2][79][20] = 1; platform_sprite[2][79][21] = 1; platform_sprite[2][79][22] = 1; platform_sprite[2][79][23] = 1; platform_sprite[2][79][24] = 1; platform_sprite[2][80][5] = 1; platform_sprite[2][80][6] = 1; platform_sprite[2][80][7] = 1; platform_sprite[2][80][8] = 1; platform_sprite[2][80][9] = 1; platform_sprite[2][80][20] = 1; platform_sprite[2][80][21] = 1; platform_sprite[2][80][22] = 1; platform_sprite[2][80][23] = 1; platform_sprite[2][80][24] = 1; platform_sprite[2][81][5] = 1; platform_sprite[2][81][6] = 1; platform_sprite[2][81][7] = 1; platform_sprite[2][81][8] = 1; platform_sprite[2][81][9] = 1; platform_sprite[2][81][20] = 1; platform_sprite[2][81][21] = 1; platform_sprite[2][81][22] = 1; platform_sprite[2][81][23] = 1; platform_sprite[2][81][24] = 1; platform_sprite[2][82][5] = 1; platform_sprite[2][82][6] = 1; platform_sprite[2][82][7] = 1; platform_sprite[2][82][8] = 1; platform_sprite[2][82][9] = 1; platform_sprite[2][82][20] = 1; platform_sprite[2][82][21] = 1; platform_sprite[2][82][22] = 1; platform_sprite[2][82][23] = 1; platform_sprite[2][82][24] = 1; platform_sprite[2][83][5] = 1; platform_sprite[2][83][6] = 1; platform_sprite[2][83][7] = 1; platform_sprite[2][83][8] = 1; platform_sprite[2][83][9] = 1; platform_sprite[2][83][20] = 1; platform_sprite[2][83][21] = 1; platform_sprite[2][83][22] = 1; platform_sprite[2][83][23] = 1; platform_sprite[2][83][24] = 1; platform_sprite[2][84][5] = 1; platform_sprite[2][84][6] = 1; platform_sprite[2][84][7] = 1; platform_sprite[2][84][8] = 1; platform_sprite[2][84][9] = 1; platform_sprite[2][84][20] = 1; platform_sprite[2][84][21] = 1; platform_sprite[2][84][22] = 1; platform_sprite[2][84][23] = 1; platform_sprite[2][84][24] = 1; platform_sprite[2][85][5] = 1; platform_sprite[2][85][6] = 1; platform_sprite[2][85][7] = 1; platform_sprite[2][85][8] = 1; platform_sprite[2][85][9] = 1; platform_sprite[2][85][20] = 1; platform_sprite[2][85][21] = 1; platform_sprite[2][85][22] = 1; platform_sprite[2][85][23] = 1; platform_sprite[2][85][24] = 1; platform_sprite[2][86][5] = 1; platform_sprite[2][86][6] = 1; platform_sprite[2][86][7] = 1; platform_sprite[2][86][8] = 1; platform_sprite[2][86][9] = 1; platform_sprite[2][86][20] = 1; platform_sprite[2][86][21] = 1; platform_sprite[2][86][22] = 1; platform_sprite[2][86][23] = 1; platform_sprite[2][86][24] = 1; platform_sprite[2][87][5] = 1; platform_sprite[2][87][6] = 1; platform_sprite[2][87][7] = 1; platform_sprite[2][87][8] = 1; platform_sprite[2][87][9] = 1; platform_sprite[2][87][20] = 1; platform_sprite[2][87][21] = 1; platform_sprite[2][87][22] = 1; platform_sprite[2][87][23] = 1; platform_sprite[2][87][24] = 1; platform_sprite[2][88][5] = 1; platform_sprite[2][88][6] = 1; platform_sprite[2][88][7] = 1; platform_sprite[2][88][8] = 1; platform_sprite[2][88][9] = 1; platform_sprite[2][88][20] = 1; platform_sprite[2][88][21] = 1; platform_sprite[2][88][22] = 1; platform_sprite[2][88][23] = 1; platform_sprite[2][88][24] = 1; platform_sprite[2][89][5] = 1; platform_sprite[2][89][6] = 1; platform_sprite[2][89][7] = 1; platform_sprite[2][89][8] = 1; platform_sprite[2][89][9] = 1; platform_sprite[2][89][20] = 1; platform_sprite[2][89][21] = 1; platform_sprite[2][89][22] = 1; platform_sprite[2][89][23] = 1; platform_sprite[2][89][24] = 1; platform_sprite[2][90][10] = 1; platform_sprite[2][90][11] = 1; platform_sprite[2][90][12] = 1; platform_sprite[2][90][13] = 1; platform_sprite[2][90][14] = 1; platform_sprite[2][90][15] = 1; platform_sprite[2][90][16] = 1; platform_sprite[2][90][17] = 1; platform_sprite[2][90][18] = 1; platform_sprite[2][90][19] = 1; platform_sprite[2][91][10] = 1; platform_sprite[2][91][11] = 1; platform_sprite[2][91][12] = 1; platform_sprite[2][91][13] = 1; platform_sprite[2][91][14] = 1; platform_sprite[2][91][15] = 1; platform_sprite[2][91][16] = 1; platform_sprite[2][91][17] = 1; platform_sprite[2][91][18] = 1; platform_sprite[2][91][19] = 1; platform_sprite[2][92][10] = 1; platform_sprite[2][92][11] = 1; platform_sprite[2][92][12] = 1; platform_sprite[2][92][13] = 1; platform_sprite[2][92][14] = 1; platform_sprite[2][92][15] = 1; platform_sprite[2][92][16] = 1; platform_sprite[2][92][17] = 1; platform_sprite[2][92][18] = 1; platform_sprite[2][92][19] = 1; platform_sprite[2][93][10] = 1; platform_sprite[2][93][11] = 1; platform_sprite[2][93][12] = 1; platform_sprite[2][93][13] = 1; platform_sprite[2][93][14] = 1; platform_sprite[2][93][15] = 1; platform_sprite[2][93][16] = 1; platform_sprite[2][93][17] = 1; platform_sprite[2][93][18] = 1; platform_sprite[2][93][19] = 1; platform_sprite[2][94][10] = 1; platform_sprite[2][94][11] = 1; platform_sprite[2][94][12] = 1; platform_sprite[2][94][13] = 1; platform_sprite[2][94][14] = 1; platform_sprite[2][94][15] = 1; platform_sprite[2][94][16] = 1; platform_sprite[2][94][17] = 1; platform_sprite[2][94][18] = 1; platform_sprite[2][94][19] = 1; 
					platform_sprite[3][5][10] = 1; platform_sprite[3][5][11] = 1; platform_sprite[3][5][12] = 1; platform_sprite[3][5][13] = 1; platform_sprite[3][5][14] = 1; platform_sprite[3][5][15] = 1; platform_sprite[3][5][16] = 1; platform_sprite[3][5][17] = 1; platform_sprite[3][5][18] = 1; platform_sprite[3][5][19] = 1; platform_sprite[3][6][10] = 1; platform_sprite[3][6][11] = 1; platform_sprite[3][6][12] = 1; platform_sprite[3][6][13] = 1; platform_sprite[3][6][14] = 1; platform_sprite[3][6][15] = 1; platform_sprite[3][6][16] = 1; platform_sprite[3][6][17] = 1; platform_sprite[3][6][18] = 1; platform_sprite[3][6][19] = 1; platform_sprite[3][7][10] = 1; platform_sprite[3][7][11] = 1; platform_sprite[3][7][12] = 1; platform_sprite[3][7][13] = 1; platform_sprite[3][7][14] = 1; platform_sprite[3][7][15] = 1; platform_sprite[3][7][16] = 1; platform_sprite[3][7][17] = 1; platform_sprite[3][7][18] = 1; platform_sprite[3][7][19] = 1; platform_sprite[3][8][10] = 1; platform_sprite[3][8][11] = 1; platform_sprite[3][8][12] = 1; platform_sprite[3][8][13] = 1; platform_sprite[3][8][14] = 1; platform_sprite[3][8][15] = 1; platform_sprite[3][8][16] = 1; platform_sprite[3][8][17] = 1; platform_sprite[3][8][18] = 1; platform_sprite[3][8][19] = 1; platform_sprite[3][9][10] = 1; platform_sprite[3][9][11] = 1; platform_sprite[3][9][12] = 1; platform_sprite[3][9][13] = 1; platform_sprite[3][9][14] = 1; platform_sprite[3][9][15] = 1; platform_sprite[3][9][16] = 1; platform_sprite[3][9][17] = 1; platform_sprite[3][9][18] = 1; platform_sprite[3][9][19] = 1; platform_sprite[3][9][20] = 1; platform_sprite[3][9][21] = 1; platform_sprite[3][9][22] = 1; platform_sprite[3][9][23] = 1; platform_sprite[3][9][24] = 1; platform_sprite[3][10][5] = 1; platform_sprite[3][10][6] = 1; platform_sprite[3][10][7] = 1; platform_sprite[3][10][8] = 1; platform_sprite[3][10][9] = 1; platform_sprite[3][10][20] = 1; platform_sprite[3][10][21] = 1; platform_sprite[3][10][22] = 1; platform_sprite[3][10][23] = 1; platform_sprite[3][10][24] = 1; platform_sprite[3][11][5] = 1; platform_sprite[3][11][6] = 1; platform_sprite[3][11][7] = 1; platform_sprite[3][11][8] = 1; platform_sprite[3][11][9] = 1; platform_sprite[3][11][20] = 1; platform_sprite[3][11][21] = 1; platform_sprite[3][11][22] = 1; platform_sprite[3][11][23] = 1; platform_sprite[3][11][24] = 1; platform_sprite[3][12][5] = 1; platform_sprite[3][12][6] = 1; platform_sprite[3][12][7] = 1; platform_sprite[3][12][8] = 1; platform_sprite[3][12][9] = 1; platform_sprite[3][12][20] = 1; platform_sprite[3][12][21] = 1; platform_sprite[3][12][22] = 1; platform_sprite[3][12][23] = 1; platform_sprite[3][12][24] = 1; platform_sprite[3][13][5] = 1; platform_sprite[3][13][6] = 1; platform_sprite[3][13][7] = 1; platform_sprite[3][13][8] = 1; platform_sprite[3][13][9] = 1; platform_sprite[3][13][20] = 1; platform_sprite[3][13][21] = 1; platform_sprite[3][13][22] = 1; platform_sprite[3][13][23] = 1; platform_sprite[3][13][24] = 1; platform_sprite[3][14][5] = 1; platform_sprite[3][14][6] = 1; platform_sprite[3][14][7] = 1; platform_sprite[3][14][8] = 1; platform_sprite[3][14][9] = 1; platform_sprite[3][14][20] = 1; platform_sprite[3][14][21] = 1; platform_sprite[3][14][22] = 1; platform_sprite[3][14][23] = 1; platform_sprite[3][14][24] = 1; platform_sprite[3][15][5] = 1; platform_sprite[3][15][6] = 1; platform_sprite[3][15][7] = 1; platform_sprite[3][15][8] = 1; platform_sprite[3][15][9] = 1; platform_sprite[3][15][20] = 1; platform_sprite[3][15][21] = 1; platform_sprite[3][15][22] = 1; platform_sprite[3][15][23] = 1; platform_sprite[3][15][24] = 1; platform_sprite[3][16][5] = 1; platform_sprite[3][16][6] = 1; platform_sprite[3][16][7] = 1; platform_sprite[3][16][8] = 1; platform_sprite[3][16][9] = 1; platform_sprite[3][16][20] = 1; platform_sprite[3][16][21] = 1; platform_sprite[3][16][22] = 1; platform_sprite[3][16][23] = 1; platform_sprite[3][16][24] = 1; platform_sprite[3][17][5] = 1; platform_sprite[3][17][6] = 1; platform_sprite[3][17][7] = 1; platform_sprite[3][17][8] = 1; platform_sprite[3][17][9] = 1; platform_sprite[3][17][20] = 1; platform_sprite[3][17][21] = 1; platform_sprite[3][17][22] = 1; platform_sprite[3][17][23] = 1; platform_sprite[3][17][24] = 1; platform_sprite[3][18][5] = 1; platform_sprite[3][18][6] = 1; platform_sprite[3][18][7] = 1; platform_sprite[3][18][8] = 1; platform_sprite[3][18][9] = 1; platform_sprite[3][18][20] = 1; platform_sprite[3][18][21] = 1; platform_sprite[3][18][22] = 1; platform_sprite[3][18][23] = 1; platform_sprite[3][18][24] = 1; platform_sprite[3][19][5] = 1; platform_sprite[3][19][6] = 1; platform_sprite[3][19][7] = 1; platform_sprite[3][19][8] = 1; platform_sprite[3][19][9] = 1; platform_sprite[3][19][20] = 1; platform_sprite[3][19][21] = 1; platform_sprite[3][19][22] = 1; platform_sprite[3][19][23] = 1; platform_sprite[3][19][24] = 1; platform_sprite[3][20][5] = 1; platform_sprite[3][20][6] = 1; platform_sprite[3][20][7] = 1; platform_sprite[3][20][8] = 1; platform_sprite[3][20][9] = 1; platform_sprite[3][20][20] = 1; platform_sprite[3][20][21] = 1; platform_sprite[3][20][22] = 1; platform_sprite[3][20][23] = 1; platform_sprite[3][20][24] = 1; platform_sprite[3][21][5] = 1; platform_sprite[3][21][6] = 1; platform_sprite[3][21][7] = 1; platform_sprite[3][21][8] = 1; platform_sprite[3][21][9] = 1; platform_sprite[3][21][20] = 1; platform_sprite[3][21][21] = 1; platform_sprite[3][21][22] = 1; platform_sprite[3][21][23] = 1; platform_sprite[3][21][24] = 1; platform_sprite[3][22][5] = 1; platform_sprite[3][22][6] = 1; platform_sprite[3][22][7] = 1; platform_sprite[3][22][8] = 1; platform_sprite[3][22][9] = 1; platform_sprite[3][22][20] = 1; platform_sprite[3][22][21] = 1; platform_sprite[3][22][22] = 1; platform_sprite[3][22][23] = 1; platform_sprite[3][22][24] = 1; platform_sprite[3][23][5] = 1; platform_sprite[3][23][6] = 1; platform_sprite[3][23][7] = 1; platform_sprite[3][23][8] = 1; platform_sprite[3][23][9] = 1; platform_sprite[3][23][20] = 1; platform_sprite[3][23][21] = 1; platform_sprite[3][23][22] = 1; platform_sprite[3][23][23] = 1; platform_sprite[3][23][24] = 1; platform_sprite[3][24][5] = 1; platform_sprite[3][24][6] = 1; platform_sprite[3][24][7] = 1; platform_sprite[3][24][8] = 1; platform_sprite[3][24][9] = 1; platform_sprite[3][24][20] = 1; platform_sprite[3][24][21] = 1; platform_sprite[3][24][22] = 1; platform_sprite[3][24][23] = 1; platform_sprite[3][24][24] = 1; platform_sprite[3][25][5] = 1; platform_sprite[3][25][6] = 1; platform_sprite[3][25][7] = 1; platform_sprite[3][25][8] = 1; platform_sprite[3][25][9] = 1; platform_sprite[3][25][20] = 1; platform_sprite[3][25][21] = 1; platform_sprite[3][25][22] = 1; platform_sprite[3][25][23] = 1; platform_sprite[3][25][24] = 1; platform_sprite[3][26][5] = 1; platform_sprite[3][26][6] = 1; platform_sprite[3][26][7] = 1; platform_sprite[3][26][8] = 1; platform_sprite[3][26][9] = 1; platform_sprite[3][26][20] = 1; platform_sprite[3][26][21] = 1; platform_sprite[3][26][22] = 1; platform_sprite[3][26][23] = 1; platform_sprite[3][26][24] = 1; platform_sprite[3][27][5] = 1; platform_sprite[3][27][6] = 1; platform_sprite[3][27][7] = 1; platform_sprite[3][27][8] = 1; platform_sprite[3][27][9] = 1; platform_sprite[3][27][20] = 1; platform_sprite[3][27][21] = 1; platform_sprite[3][27][22] = 1; platform_sprite[3][27][23] = 1; platform_sprite[3][27][24] = 1; platform_sprite[3][28][5] = 1; platform_sprite[3][28][6] = 1; platform_sprite[3][28][7] = 1; platform_sprite[3][28][8] = 1; platform_sprite[3][28][9] = 1; platform_sprite[3][28][20] = 1; platform_sprite[3][28][21] = 1; platform_sprite[3][28][22] = 1; platform_sprite[3][28][23] = 1; platform_sprite[3][28][24] = 1; platform_sprite[3][29][5] = 1; platform_sprite[3][29][6] = 1; platform_sprite[3][29][7] = 1; platform_sprite[3][29][8] = 1; platform_sprite[3][29][9] = 1; platform_sprite[3][29][20] = 1; platform_sprite[3][29][21] = 1; platform_sprite[3][29][22] = 1; platform_sprite[3][29][23] = 1; platform_sprite[3][29][24] = 1; platform_sprite[3][30][5] = 1; platform_sprite[3][30][6] = 1; platform_sprite[3][30][7] = 1; platform_sprite[3][30][8] = 1; platform_sprite[3][30][9] = 1; platform_sprite[3][30][20] = 1; platform_sprite[3][30][21] = 1; platform_sprite[3][30][22] = 1; platform_sprite[3][30][23] = 1; platform_sprite[3][30][24] = 1; platform_sprite[3][31][5] = 1; platform_sprite[3][31][6] = 1; platform_sprite[3][31][7] = 1; platform_sprite[3][31][8] = 1; platform_sprite[3][31][9] = 1; platform_sprite[3][31][20] = 1; platform_sprite[3][31][21] = 1; platform_sprite[3][31][22] = 1; platform_sprite[3][31][23] = 1; platform_sprite[3][31][24] = 1; platform_sprite[3][32][5] = 1; platform_sprite[3][32][6] = 1; platform_sprite[3][32][7] = 1; platform_sprite[3][32][8] = 1; platform_sprite[3][32][9] = 1; platform_sprite[3][32][20] = 1; platform_sprite[3][32][21] = 1; platform_sprite[3][32][22] = 1; platform_sprite[3][32][23] = 1; platform_sprite[3][32][24] = 1; platform_sprite[3][33][5] = 1; platform_sprite[3][33][6] = 1; platform_sprite[3][33][7] = 1; platform_sprite[3][33][8] = 1; platform_sprite[3][33][9] = 1; platform_sprite[3][33][20] = 1; platform_sprite[3][33][21] = 1; platform_sprite[3][33][22] = 1; platform_sprite[3][33][23] = 1; platform_sprite[3][33][24] = 1; platform_sprite[3][34][5] = 1; platform_sprite[3][34][6] = 1; platform_sprite[3][34][7] = 1; platform_sprite[3][34][8] = 1; platform_sprite[3][34][9] = 1; platform_sprite[3][34][20] = 1; platform_sprite[3][34][21] = 1; platform_sprite[3][34][22] = 1; platform_sprite[3][34][23] = 1; platform_sprite[3][34][24] = 1; platform_sprite[3][35][5] = 1; platform_sprite[3][35][6] = 1; platform_sprite[3][35][7] = 1; platform_sprite[3][35][8] = 1; platform_sprite[3][35][9] = 1; platform_sprite[3][35][20] = 1; platform_sprite[3][35][21] = 1; platform_sprite[3][35][22] = 1; platform_sprite[3][35][23] = 1; platform_sprite[3][35][24] = 1; platform_sprite[3][36][5] = 1; platform_sprite[3][36][6] = 1; platform_sprite[3][36][7] = 1; platform_sprite[3][36][8] = 1; platform_sprite[3][36][9] = 1; platform_sprite[3][36][20] = 1; platform_sprite[3][36][21] = 1; platform_sprite[3][36][22] = 1; platform_sprite[3][36][23] = 1; platform_sprite[3][36][24] = 1; platform_sprite[3][37][5] = 1; platform_sprite[3][37][6] = 1; platform_sprite[3][37][7] = 1; platform_sprite[3][37][8] = 1; platform_sprite[3][37][9] = 1; platform_sprite[3][37][20] = 1; platform_sprite[3][37][21] = 1; platform_sprite[3][37][22] = 1; platform_sprite[3][37][23] = 1; platform_sprite[3][37][24] = 1; platform_sprite[3][38][5] = 1; platform_sprite[3][38][6] = 1; platform_sprite[3][38][7] = 1; platform_sprite[3][38][8] = 1; platform_sprite[3][38][9] = 1; platform_sprite[3][38][20] = 1; platform_sprite[3][38][21] = 1; platform_sprite[3][38][22] = 1; platform_sprite[3][38][23] = 1; platform_sprite[3][38][24] = 1; platform_sprite[3][39][5] = 1; platform_sprite[3][39][6] = 1; platform_sprite[3][39][7] = 1; platform_sprite[3][39][8] = 1; platform_sprite[3][39][9] = 1; platform_sprite[3][39][20] = 1; platform_sprite[3][39][21] = 1; platform_sprite[3][39][22] = 1; platform_sprite[3][39][23] = 1; platform_sprite[3][39][24] = 1; platform_sprite[3][40][5] = 1; platform_sprite[3][40][6] = 1; platform_sprite[3][40][7] = 1; platform_sprite[3][40][8] = 1; platform_sprite[3][40][9] = 1; platform_sprite[3][40][20] = 1; platform_sprite[3][40][21] = 1; platform_sprite[3][40][22] = 1; platform_sprite[3][40][23] = 1; platform_sprite[3][40][24] = 1; platform_sprite[3][41][5] = 1; platform_sprite[3][41][6] = 1; platform_sprite[3][41][7] = 1; platform_sprite[3][41][8] = 1; platform_sprite[3][41][9] = 1; platform_sprite[3][41][20] = 1; platform_sprite[3][41][21] = 1; platform_sprite[3][41][22] = 1; platform_sprite[3][41][23] = 1; platform_sprite[3][41][24] = 1; platform_sprite[3][42][5] = 1; platform_sprite[3][42][6] = 1; platform_sprite[3][42][7] = 1; platform_sprite[3][42][8] = 1; platform_sprite[3][42][9] = 1; platform_sprite[3][42][20] = 1; platform_sprite[3][42][21] = 1; platform_sprite[3][42][22] = 1; platform_sprite[3][42][23] = 1; platform_sprite[3][42][24] = 1; platform_sprite[3][43][5] = 1; platform_sprite[3][43][6] = 1; platform_sprite[3][43][7] = 1; platform_sprite[3][43][8] = 1; platform_sprite[3][43][9] = 1; platform_sprite[3][43][20] = 1; platform_sprite[3][43][21] = 1; platform_sprite[3][43][22] = 1; platform_sprite[3][43][23] = 1; platform_sprite[3][43][24] = 1; platform_sprite[3][44][5] = 1; platform_sprite[3][44][6] = 1; platform_sprite[3][44][7] = 1; platform_sprite[3][44][8] = 1; platform_sprite[3][44][9] = 1; platform_sprite[3][44][20] = 1; platform_sprite[3][44][21] = 1; platform_sprite[3][44][22] = 1; platform_sprite[3][44][23] = 1; platform_sprite[3][44][24] = 1; platform_sprite[3][45][5] = 1; platform_sprite[3][45][6] = 1; platform_sprite[3][45][7] = 1; platform_sprite[3][45][8] = 1; platform_sprite[3][45][9] = 1; platform_sprite[3][45][20] = 1; platform_sprite[3][45][21] = 1; platform_sprite[3][45][22] = 1; platform_sprite[3][45][23] = 1; platform_sprite[3][45][24] = 1; platform_sprite[3][46][5] = 1; platform_sprite[3][46][6] = 1; platform_sprite[3][46][7] = 1; platform_sprite[3][46][8] = 1; platform_sprite[3][46][9] = 1; platform_sprite[3][46][20] = 1; platform_sprite[3][46][21] = 1; platform_sprite[3][46][22] = 1; platform_sprite[3][46][23] = 1; platform_sprite[3][46][24] = 1; platform_sprite[3][47][5] = 1; platform_sprite[3][47][6] = 1; platform_sprite[3][47][7] = 1; platform_sprite[3][47][8] = 1; platform_sprite[3][47][9] = 1; platform_sprite[3][47][20] = 1; platform_sprite[3][47][21] = 1; platform_sprite[3][47][22] = 1; platform_sprite[3][47][23] = 1; platform_sprite[3][47][24] = 1; platform_sprite[3][48][5] = 1; platform_sprite[3][48][6] = 1; platform_sprite[3][48][7] = 1; platform_sprite[3][48][8] = 1; platform_sprite[3][48][9] = 1; platform_sprite[3][48][20] = 1; platform_sprite[3][48][21] = 1; platform_sprite[3][48][22] = 1; platform_sprite[3][48][23] = 1; platform_sprite[3][48][24] = 1; platform_sprite[3][49][5] = 1; platform_sprite[3][49][6] = 1; platform_sprite[3][49][7] = 1; platform_sprite[3][49][8] = 1; platform_sprite[3][49][9] = 1; platform_sprite[3][49][20] = 1; platform_sprite[3][49][21] = 1; platform_sprite[3][49][22] = 1; platform_sprite[3][49][23] = 1; platform_sprite[3][49][24] = 1; platform_sprite[3][50][5] = 1; platform_sprite[3][50][6] = 1; platform_sprite[3][50][7] = 1; platform_sprite[3][50][8] = 1; platform_sprite[3][50][9] = 1; platform_sprite[3][50][20] = 1; platform_sprite[3][50][21] = 1; platform_sprite[3][50][22] = 1; platform_sprite[3][50][23] = 1; platform_sprite[3][50][24] = 1; platform_sprite[3][51][5] = 1; platform_sprite[3][51][6] = 1; platform_sprite[3][51][7] = 1; platform_sprite[3][51][8] = 1; platform_sprite[3][51][9] = 1; platform_sprite[3][51][20] = 1; platform_sprite[3][51][21] = 1; platform_sprite[3][51][22] = 1; platform_sprite[3][51][23] = 1; platform_sprite[3][51][24] = 1; platform_sprite[3][52][5] = 1; platform_sprite[3][52][6] = 1; platform_sprite[3][52][7] = 1; platform_sprite[3][52][8] = 1; platform_sprite[3][52][9] = 1; platform_sprite[3][52][20] = 1; platform_sprite[3][52][21] = 1; platform_sprite[3][52][22] = 1; platform_sprite[3][52][23] = 1; platform_sprite[3][52][24] = 1; platform_sprite[3][53][5] = 1; platform_sprite[3][53][6] = 1; platform_sprite[3][53][7] = 1; platform_sprite[3][53][8] = 1; platform_sprite[3][53][9] = 1; platform_sprite[3][53][20] = 1; platform_sprite[3][53][21] = 1; platform_sprite[3][53][22] = 1; platform_sprite[3][53][23] = 1; platform_sprite[3][53][24] = 1; platform_sprite[3][54][5] = 1; platform_sprite[3][54][6] = 1; platform_sprite[3][54][7] = 1; platform_sprite[3][54][8] = 1; platform_sprite[3][54][9] = 1; platform_sprite[3][54][20] = 1; platform_sprite[3][54][21] = 1; platform_sprite[3][54][22] = 1; platform_sprite[3][54][23] = 1; platform_sprite[3][54][24] = 1; platform_sprite[3][55][5] = 1; platform_sprite[3][55][6] = 1; platform_sprite[3][55][7] = 1; platform_sprite[3][55][8] = 1; platform_sprite[3][55][9] = 1; platform_sprite[3][55][20] = 1; platform_sprite[3][55][21] = 1; platform_sprite[3][55][22] = 1; platform_sprite[3][55][23] = 1; platform_sprite[3][55][24] = 1; platform_sprite[3][56][5] = 1; platform_sprite[3][56][6] = 1; platform_sprite[3][56][7] = 1; platform_sprite[3][56][8] = 1; platform_sprite[3][56][9] = 1; platform_sprite[3][56][20] = 1; platform_sprite[3][56][21] = 1; platform_sprite[3][56][22] = 1; platform_sprite[3][56][23] = 1; platform_sprite[3][56][24] = 1; platform_sprite[3][57][5] = 1; platform_sprite[3][57][6] = 1; platform_sprite[3][57][7] = 1; platform_sprite[3][57][8] = 1; platform_sprite[3][57][9] = 1; platform_sprite[3][57][20] = 1; platform_sprite[3][57][21] = 1; platform_sprite[3][57][22] = 1; platform_sprite[3][57][23] = 1; platform_sprite[3][57][24] = 1; platform_sprite[3][58][5] = 1; platform_sprite[3][58][6] = 1; platform_sprite[3][58][7] = 1; platform_sprite[3][58][8] = 1; platform_sprite[3][58][9] = 1; platform_sprite[3][58][20] = 1; platform_sprite[3][58][21] = 1; platform_sprite[3][58][22] = 1; platform_sprite[3][58][23] = 1; platform_sprite[3][58][24] = 1; platform_sprite[3][59][5] = 1; platform_sprite[3][59][6] = 1; platform_sprite[3][59][7] = 1; platform_sprite[3][59][8] = 1; platform_sprite[3][59][9] = 1; platform_sprite[3][59][20] = 1; platform_sprite[3][59][21] = 1; platform_sprite[3][59][22] = 1; platform_sprite[3][59][23] = 1; platform_sprite[3][59][24] = 1; platform_sprite[3][60][5] = 1; platform_sprite[3][60][6] = 1; platform_sprite[3][60][7] = 1; platform_sprite[3][60][8] = 1; platform_sprite[3][60][9] = 1; platform_sprite[3][60][20] = 1; platform_sprite[3][60][21] = 1; platform_sprite[3][60][22] = 1; platform_sprite[3][60][23] = 1; platform_sprite[3][60][24] = 1; platform_sprite[3][61][5] = 1; platform_sprite[3][61][6] = 1; platform_sprite[3][61][7] = 1; platform_sprite[3][61][8] = 1; platform_sprite[3][61][9] = 1; platform_sprite[3][61][20] = 1; platform_sprite[3][61][21] = 1; platform_sprite[3][61][22] = 1; platform_sprite[3][61][23] = 1; platform_sprite[3][61][24] = 1; platform_sprite[3][62][5] = 1; platform_sprite[3][62][6] = 1; platform_sprite[3][62][7] = 1; platform_sprite[3][62][8] = 1; platform_sprite[3][62][9] = 1; platform_sprite[3][62][20] = 1; platform_sprite[3][62][21] = 1; platform_sprite[3][62][22] = 1; platform_sprite[3][62][23] = 1; platform_sprite[3][62][24] = 1; platform_sprite[3][63][5] = 1; platform_sprite[3][63][6] = 1; platform_sprite[3][63][7] = 1; platform_sprite[3][63][8] = 1; platform_sprite[3][63][9] = 1; platform_sprite[3][63][20] = 1; platform_sprite[3][63][21] = 1; platform_sprite[3][63][22] = 1; platform_sprite[3][63][23] = 1; platform_sprite[3][63][24] = 1; platform_sprite[3][64][5] = 1; platform_sprite[3][64][6] = 1; platform_sprite[3][64][7] = 1; platform_sprite[3][64][8] = 1; platform_sprite[3][64][9] = 1; platform_sprite[3][64][20] = 1; platform_sprite[3][64][21] = 1; platform_sprite[3][64][22] = 1; platform_sprite[3][64][23] = 1; platform_sprite[3][64][24] = 1; platform_sprite[3][65][5] = 1; platform_sprite[3][65][6] = 1; platform_sprite[3][65][7] = 1; platform_sprite[3][65][8] = 1; platform_sprite[3][65][9] = 1; platform_sprite[3][65][20] = 1; platform_sprite[3][65][21] = 1; platform_sprite[3][65][22] = 1; platform_sprite[3][65][23] = 1; platform_sprite[3][65][24] = 1; platform_sprite[3][66][5] = 1; platform_sprite[3][66][6] = 1; platform_sprite[3][66][7] = 1; platform_sprite[3][66][8] = 1; platform_sprite[3][66][9] = 1; platform_sprite[3][66][20] = 1; platform_sprite[3][66][21] = 1; platform_sprite[3][66][22] = 1; platform_sprite[3][66][23] = 1; platform_sprite[3][66][24] = 1; platform_sprite[3][67][5] = 1; platform_sprite[3][67][6] = 1; platform_sprite[3][67][7] = 1; platform_sprite[3][67][8] = 1; platform_sprite[3][67][9] = 1; platform_sprite[3][67][20] = 1; platform_sprite[3][67][21] = 1; platform_sprite[3][67][22] = 1; platform_sprite[3][67][23] = 1; platform_sprite[3][67][24] = 1; platform_sprite[3][68][5] = 1; platform_sprite[3][68][6] = 1; platform_sprite[3][68][7] = 1; platform_sprite[3][68][8] = 1; platform_sprite[3][68][9] = 1; platform_sprite[3][68][20] = 1; platform_sprite[3][68][21] = 1; platform_sprite[3][68][22] = 1; platform_sprite[3][68][23] = 1; platform_sprite[3][68][24] = 1; platform_sprite[3][69][5] = 1; platform_sprite[3][69][6] = 1; platform_sprite[3][69][7] = 1; platform_sprite[3][69][8] = 1; platform_sprite[3][69][9] = 1; platform_sprite[3][69][20] = 1; platform_sprite[3][69][21] = 1; platform_sprite[3][69][22] = 1; platform_sprite[3][69][23] = 1; platform_sprite[3][69][24] = 1; platform_sprite[3][70][5] = 1; platform_sprite[3][70][6] = 1; platform_sprite[3][70][7] = 1; platform_sprite[3][70][8] = 1; platform_sprite[3][70][9] = 1; platform_sprite[3][70][20] = 1; platform_sprite[3][70][21] = 1; platform_sprite[3][70][22] = 1; platform_sprite[3][70][23] = 1; platform_sprite[3][70][24] = 1; platform_sprite[3][71][5] = 1; platform_sprite[3][71][6] = 1; platform_sprite[3][71][7] = 1; platform_sprite[3][71][8] = 1; platform_sprite[3][71][9] = 1; platform_sprite[3][71][20] = 1; platform_sprite[3][71][21] = 1; platform_sprite[3][71][22] = 1; platform_sprite[3][71][23] = 1; platform_sprite[3][71][24] = 1; platform_sprite[3][72][5] = 1; platform_sprite[3][72][6] = 1; platform_sprite[3][72][7] = 1; platform_sprite[3][72][8] = 1; platform_sprite[3][72][9] = 1; platform_sprite[3][72][20] = 1; platform_sprite[3][72][21] = 1; platform_sprite[3][72][22] = 1; platform_sprite[3][72][23] = 1; platform_sprite[3][72][24] = 1; platform_sprite[3][73][5] = 1; platform_sprite[3][73][6] = 1; platform_sprite[3][73][7] = 1; platform_sprite[3][73][8] = 1; platform_sprite[3][73][9] = 1; platform_sprite[3][73][20] = 1; platform_sprite[3][73][21] = 1; platform_sprite[3][73][22] = 1; platform_sprite[3][73][23] = 1; platform_sprite[3][73][24] = 1; platform_sprite[3][74][5] = 1; platform_sprite[3][74][6] = 1; platform_sprite[3][74][7] = 1; platform_sprite[3][74][8] = 1; platform_sprite[3][74][9] = 1; platform_sprite[3][74][20] = 1; platform_sprite[3][74][21] = 1; platform_sprite[3][74][22] = 1; platform_sprite[3][74][23] = 1; platform_sprite[3][74][24] = 1; platform_sprite[3][75][5] = 1; platform_sprite[3][75][6] = 1; platform_sprite[3][75][7] = 1; platform_sprite[3][75][8] = 1; platform_sprite[3][75][9] = 1; platform_sprite[3][75][20] = 1; platform_sprite[3][75][21] = 1; platform_sprite[3][75][22] = 1; platform_sprite[3][75][23] = 1; platform_sprite[3][75][24] = 1; platform_sprite[3][76][5] = 1; platform_sprite[3][76][6] = 1; platform_sprite[3][76][7] = 1; platform_sprite[3][76][8] = 1; platform_sprite[3][76][9] = 1; platform_sprite[3][76][20] = 1; platform_sprite[3][76][21] = 1; platform_sprite[3][76][22] = 1; platform_sprite[3][76][23] = 1; platform_sprite[3][76][24] = 1; platform_sprite[3][77][5] = 1; platform_sprite[3][77][6] = 1; platform_sprite[3][77][7] = 1; platform_sprite[3][77][8] = 1; platform_sprite[3][77][9] = 1; platform_sprite[3][77][20] = 1; platform_sprite[3][77][21] = 1; platform_sprite[3][77][22] = 1; platform_sprite[3][77][23] = 1; platform_sprite[3][77][24] = 1; platform_sprite[3][78][5] = 1; platform_sprite[3][78][6] = 1; platform_sprite[3][78][7] = 1; platform_sprite[3][78][8] = 1; platform_sprite[3][78][9] = 1; platform_sprite[3][78][20] = 1; platform_sprite[3][78][21] = 1; platform_sprite[3][78][22] = 1; platform_sprite[3][78][23] = 1; platform_sprite[3][78][24] = 1; platform_sprite[3][79][5] = 1; platform_sprite[3][79][6] = 1; platform_sprite[3][79][7] = 1; platform_sprite[3][79][8] = 1; platform_sprite[3][79][9] = 1; platform_sprite[3][79][20] = 1; platform_sprite[3][79][21] = 1; platform_sprite[3][79][22] = 1; platform_sprite[3][79][23] = 1; platform_sprite[3][79][24] = 1; platform_sprite[3][80][5] = 1; platform_sprite[3][80][6] = 1; platform_sprite[3][80][7] = 1; platform_sprite[3][80][8] = 1; platform_sprite[3][80][9] = 1; platform_sprite[3][80][20] = 1; platform_sprite[3][80][21] = 1; platform_sprite[3][80][22] = 1; platform_sprite[3][80][23] = 1; platform_sprite[3][80][24] = 1; platform_sprite[3][81][5] = 1; platform_sprite[3][81][6] = 1; platform_sprite[3][81][7] = 1; platform_sprite[3][81][8] = 1; platform_sprite[3][81][9] = 1; platform_sprite[3][81][20] = 1; platform_sprite[3][81][21] = 1; platform_sprite[3][81][22] = 1; platform_sprite[3][81][23] = 1; platform_sprite[3][81][24] = 1; platform_sprite[3][82][5] = 1; platform_sprite[3][82][6] = 1; platform_sprite[3][82][7] = 1; platform_sprite[3][82][8] = 1; platform_sprite[3][82][9] = 1; platform_sprite[3][82][20] = 1; platform_sprite[3][82][21] = 1; platform_sprite[3][82][22] = 1; platform_sprite[3][82][23] = 1; platform_sprite[3][82][24] = 1; platform_sprite[3][83][5] = 1; platform_sprite[3][83][6] = 1; platform_sprite[3][83][7] = 1; platform_sprite[3][83][8] = 1; platform_sprite[3][83][9] = 1; platform_sprite[3][83][20] = 1; platform_sprite[3][83][21] = 1; platform_sprite[3][83][22] = 1; platform_sprite[3][83][23] = 1; platform_sprite[3][83][24] = 1; platform_sprite[3][84][5] = 1; platform_sprite[3][84][6] = 1; platform_sprite[3][84][7] = 1; platform_sprite[3][84][8] = 1; platform_sprite[3][84][9] = 1; platform_sprite[3][84][20] = 1; platform_sprite[3][84][21] = 1; platform_sprite[3][84][22] = 1; platform_sprite[3][84][23] = 1; platform_sprite[3][84][24] = 1; platform_sprite[3][85][5] = 1; platform_sprite[3][85][6] = 1; platform_sprite[3][85][7] = 1; platform_sprite[3][85][8] = 1; platform_sprite[3][85][9] = 1; platform_sprite[3][85][20] = 1; platform_sprite[3][85][21] = 1; platform_sprite[3][85][22] = 1; platform_sprite[3][85][23] = 1; platform_sprite[3][85][24] = 1; platform_sprite[3][86][5] = 1; platform_sprite[3][86][6] = 1; platform_sprite[3][86][7] = 1; platform_sprite[3][86][8] = 1; platform_sprite[3][86][9] = 1; platform_sprite[3][86][20] = 1; platform_sprite[3][86][21] = 1; platform_sprite[3][86][22] = 1; platform_sprite[3][86][23] = 1; platform_sprite[3][86][24] = 1; platform_sprite[3][87][5] = 1; platform_sprite[3][87][6] = 1; platform_sprite[3][87][7] = 1; platform_sprite[3][87][8] = 1; platform_sprite[3][87][9] = 1; platform_sprite[3][87][20] = 1; platform_sprite[3][87][21] = 1; platform_sprite[3][87][22] = 1; platform_sprite[3][87][23] = 1; platform_sprite[3][87][24] = 1; platform_sprite[3][88][5] = 1; platform_sprite[3][88][6] = 1; platform_sprite[3][88][7] = 1; platform_sprite[3][88][8] = 1; platform_sprite[3][88][9] = 1; platform_sprite[3][88][20] = 1; platform_sprite[3][88][21] = 1; platform_sprite[3][88][22] = 1; platform_sprite[3][88][23] = 1; platform_sprite[3][88][24] = 1; platform_sprite[3][89][5] = 1; platform_sprite[3][89][6] = 1; platform_sprite[3][89][7] = 1; platform_sprite[3][89][8] = 1; platform_sprite[3][89][9] = 1; platform_sprite[3][89][20] = 1; platform_sprite[3][89][21] = 1; platform_sprite[3][89][22] = 1; platform_sprite[3][89][23] = 1; platform_sprite[3][89][24] = 1; platform_sprite[3][90][10] = 1; platform_sprite[3][90][11] = 1; platform_sprite[3][90][12] = 1; platform_sprite[3][90][13] = 1; platform_sprite[3][90][14] = 1; platform_sprite[3][90][15] = 1; platform_sprite[3][90][16] = 1; platform_sprite[3][90][17] = 1; platform_sprite[3][90][18] = 1; platform_sprite[3][90][19] = 1; platform_sprite[3][91][10] = 1; platform_sprite[3][91][11] = 1; platform_sprite[3][91][12] = 1; platform_sprite[3][91][13] = 1; platform_sprite[3][91][14] = 1; platform_sprite[3][91][15] = 1; platform_sprite[3][91][16] = 1; platform_sprite[3][91][17] = 1; platform_sprite[3][91][18] = 1; platform_sprite[3][91][19] = 1; platform_sprite[3][92][10] = 1; platform_sprite[3][92][11] = 1; platform_sprite[3][92][12] = 1; platform_sprite[3][92][13] = 1; platform_sprite[3][92][14] = 1; platform_sprite[3][92][15] = 1; platform_sprite[3][92][16] = 1; platform_sprite[3][92][17] = 1; platform_sprite[3][92][18] = 1; platform_sprite[3][92][19] = 1; platform_sprite[3][93][10] = 1; platform_sprite[3][93][11] = 1; platform_sprite[3][93][12] = 1; platform_sprite[3][93][13] = 1; platform_sprite[3][93][14] = 1; platform_sprite[3][93][15] = 1; platform_sprite[3][93][16] = 1; platform_sprite[3][93][17] = 1; platform_sprite[3][93][18] = 1; platform_sprite[3][93][19] = 1; platform_sprite[3][94][10] = 1; platform_sprite[3][94][11] = 1; platform_sprite[3][94][12] = 1; platform_sprite[3][94][13] = 1; platform_sprite[3][94][14] = 1; platform_sprite[3][94][15] = 1; platform_sprite[3][94][16] = 1; platform_sprite[3][94][17] = 1; platform_sprite[3][94][18] = 1; platform_sprite[3][94][19] = 1; 
						
					//platform painting
					for (i = 0; i < 4; i = i + 1) begin
						if (platform_v[i] >= 0 && platform_v[i] <= 30 && platform_h[i] >= 0 && platform_h[i] <= 100) begin
							if (platform_sprite[i][platform_h[i]][platform_v[i]] == 1) begin
								r = 0;
								g = 0;
								b = 0;
							end
						end
					end
					//----------------------------------
					
					//doodle painting----------------------
					if (doodle_v >= 0 && doodle_v <= 80 && doodle_h >= 0 && doodle_h <= 80) begin
						if (doodle_sprite[sprite_choice][doodle_h][doodle_v] == 1) begin
							r = 0;
							g = 0;
							b = 0;
						end
						else if (doodle_sprite[sprite_choice][doodle_h][doodle_v] == 2) begin
							r = 0;
							g = 1;
							b = 0;
						end
					end
					
					//drawing the frame
					if (((count_v <= 5  || count_v >= 760) && count_h >= 342 && count_h <= 682) || (count_h >= 342 && count_h <= 346) || (count_h >= 677 && count_h <= 682)) begin
							r = 0;
							g = 0;
							b = 0;
						end
					//---
				end
				//if the game is over---
				else 
					begin
					//background painting
					if (count_h >= 0) 
						begin
						r = 0;
						g = 0;
						b = 0;
						end
					//drawing the frame
					if (((count_v <= 5  || count_v >= 760) && count_h >= 342 && count_h <= 682) || (count_h >= 342 && count_h <= 346) || (count_h >= 677 && count_h <= 682))
						begin
						r = 1;
						g = 1;
						b = 1;
						end
					//---
					end
				end //EA ends
				
			//out of screen---------
			else begin
				r = 0;
				g = 0;
				b = 0;
			end
			//---------------------
			
	end
endmodule